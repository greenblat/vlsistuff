`celldefine
module BUF (input A, output Y);
assign  Y = A;
endmodule
`endcelldefine
