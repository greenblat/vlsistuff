
`timescale 1ns/1ps
module tb;
parameter IDWID=4; parameter DWID=64; parameter EXTRAS=8; parameter WSTRB=DWID/8;

reg [31:0] cycles;   initial cycles=0;
reg [31:0] errors;   initial errors=0;
reg [31:0] wrongs;   initial wrongs=0;
reg [31:0] Panics;   initial Panics=0;
reg [31:0] corrects; initial corrects=0;
reg [31:0] marker;   initial marker=0;
reg [31:0] marker0;   initial marker0=0;
reg [31:0] marker1;   initial marker1=0;
reg [31:0] marker2;   initial marker2=0;
reg [31:0] marker3;   initial marker3=0;
reg [31:0] Index;   initial Index=0;



reg clk; reg rst_n;
always begin
    clk = 0;
    #10;
    clk = 1;
    #3;
    $python("negedge()");
    #3;
    $python("auxs()");
    #4;
end
initial begin
    $dumpvars(0,tb);
    rst_n = 0;
    #100;
    rst_n = 1;
end

reg  [2:0] slv0_awsize ; initial slv0_awsize = 0;
reg  [2:0] slv0_arsize ; initial slv0_arsize = 0;

wire  [IDWID-1:0] slv0_arid ;
wire  [31:0] slv0_araddr ;
wire  [7:0] slv0_arlen ;
wire  [EXTRAS-1:0] slv0_arextras ;
wire  [1:0] slv0_arburst ;
wire  slv0_arvalid ;
reg  slv0_arready ;
reg  [IDWID-1:0] slv0_rid ;
reg  [DWID-1:0] slv0_rdata ;
reg  [1:0] slv0_rresp ;
reg  slv0_rlast ;
reg  slv0_rvalid ;
wire  slv0_rready ;

wire  [IDWID-1:0] slv0_awid ;
wire  [31:0] slv0_awaddr ;
wire  [7:0] slv0_awlen ;
wire  [EXTRAS-1:0] slv0_awextras ;
wire  [1:0] slv0_awburst ;
wire  slv0_awvalid ;
reg  slv0_awready ;
wire  [DWID-1:0] slv0_wdata ;
wire  [WSTRB-1:0] slv0_wstrb ;
wire  slv0_wlast ;
wire  slv0_wvalid ;
reg  slv0_wready ;
reg  [IDWID-1:0] slv0_bid ;
reg  [1:0] slv0_bresp ;
reg  slv0_bvalid ;
wire  slv0_bready ;

initial slv0_arready = 0;
initial slv0_awready = 0;
initial slv0_rvalid = 0;
initial slv0_bvalid = 0;

reg  [2:0] slv1_awsize ; initial slv1_awsize = 0;
reg  [2:0] slv1_arsize ; initial slv1_arsize = 0;

wire  [IDWID-1:0] slv1_arid ;
wire  [31:0] slv1_araddr ;
wire  [7:0] slv1_arlen ;
wire  [EXTRAS-1:0] slv1_arextras ;
wire  [1:0] slv1_arburst ;
wire  slv1_arvalid ;
reg  slv1_arready ;
reg  [IDWID-1:0] slv1_rid ;
reg  [DWID-1:0] slv1_rdata ;
reg  [1:0] slv1_rresp ;
reg  slv1_rlast ;
reg  slv1_rvalid ;
wire  slv1_rready ;

wire  [IDWID-1:0] slv1_awid ;
wire  [31:0] slv1_awaddr ;
wire  [7:0] slv1_awlen ;
wire  [EXTRAS-1:0] slv1_awextras ;
wire  [1:0] slv1_awburst ;
wire  slv1_awvalid ;
reg  slv1_awready ;
wire  [DWID-1:0] slv1_wdata ;
wire  [WSTRB-1:0] slv1_wstrb ;
wire  slv1_wlast ;
wire  slv1_wvalid ;
reg  slv1_wready ;
reg  [IDWID-1:0] slv1_bid ;
reg  [1:0] slv1_bresp ;
reg  slv1_bvalid ;
wire  slv1_bready ;

initial slv1_arready = 0;
initial slv1_awready = 0;
initial slv1_rvalid = 0;
initial slv1_bvalid = 0;

reg  [2:0] slv10_awsize ; initial slv10_awsize = 0;
reg  [2:0] slv10_arsize ; initial slv10_arsize = 0;

wire  [IDWID-1:0] slv10_arid ;
wire  [31:0] slv10_araddr ;
wire  [7:0] slv10_arlen ;
wire  [EXTRAS-1:0] slv10_arextras ;
wire  [1:0] slv10_arburst ;
wire  slv10_arvalid ;
reg  slv10_arready ;
reg  [IDWID-1:0] slv10_rid ;
reg  [DWID-1:0] slv10_rdata ;
reg  [1:0] slv10_rresp ;
reg  slv10_rlast ;
reg  slv10_rvalid ;
wire  slv10_rready ;

wire  [IDWID-1:0] slv10_awid ;
wire  [31:0] slv10_awaddr ;
wire  [7:0] slv10_awlen ;
wire  [EXTRAS-1:0] slv10_awextras ;
wire  [1:0] slv10_awburst ;
wire  slv10_awvalid ;
reg  slv10_awready ;
wire  [DWID-1:0] slv10_wdata ;
wire  [WSTRB-1:0] slv10_wstrb ;
wire  slv10_wlast ;
wire  slv10_wvalid ;
reg  slv10_wready ;
reg  [IDWID-1:0] slv10_bid ;
reg  [1:0] slv10_bresp ;
reg  slv10_bvalid ;
wire  slv10_bready ;

initial slv10_arready = 0;
initial slv10_awready = 0;
initial slv10_rvalid = 0;
initial slv10_bvalid = 0;

reg  [2:0] slv11_awsize ; initial slv11_awsize = 0;
reg  [2:0] slv11_arsize ; initial slv11_arsize = 0;

wire  [IDWID-1:0] slv11_arid ;
wire  [31:0] slv11_araddr ;
wire  [7:0] slv11_arlen ;
wire  [EXTRAS-1:0] slv11_arextras ;
wire  [1:0] slv11_arburst ;
wire  slv11_arvalid ;
reg  slv11_arready ;
reg  [IDWID-1:0] slv11_rid ;
reg  [DWID-1:0] slv11_rdata ;
reg  [1:0] slv11_rresp ;
reg  slv11_rlast ;
reg  slv11_rvalid ;
wire  slv11_rready ;

wire  [IDWID-1:0] slv11_awid ;
wire  [31:0] slv11_awaddr ;
wire  [7:0] slv11_awlen ;
wire  [EXTRAS-1:0] slv11_awextras ;
wire  [1:0] slv11_awburst ;
wire  slv11_awvalid ;
reg  slv11_awready ;
wire  [DWID-1:0] slv11_wdata ;
wire  [WSTRB-1:0] slv11_wstrb ;
wire  slv11_wlast ;
wire  slv11_wvalid ;
reg  slv11_wready ;
reg  [IDWID-1:0] slv11_bid ;
reg  [1:0] slv11_bresp ;
reg  slv11_bvalid ;
wire  slv11_bready ;

initial slv11_arready = 0;
initial slv11_awready = 0;
initial slv11_rvalid = 0;
initial slv11_bvalid = 0;

reg  [2:0] slv12_awsize ; initial slv12_awsize = 0;
reg  [2:0] slv12_arsize ; initial slv12_arsize = 0;

wire  [IDWID-1:0] slv12_arid ;
wire  [31:0] slv12_araddr ;
wire  [7:0] slv12_arlen ;
wire  [EXTRAS-1:0] slv12_arextras ;
wire  [1:0] slv12_arburst ;
wire  slv12_arvalid ;
reg  slv12_arready ;
reg  [IDWID-1:0] slv12_rid ;
reg  [DWID-1:0] slv12_rdata ;
reg  [1:0] slv12_rresp ;
reg  slv12_rlast ;
reg  slv12_rvalid ;
wire  slv12_rready ;

wire  [IDWID-1:0] slv12_awid ;
wire  [31:0] slv12_awaddr ;
wire  [7:0] slv12_awlen ;
wire  [EXTRAS-1:0] slv12_awextras ;
wire  [1:0] slv12_awburst ;
wire  slv12_awvalid ;
reg  slv12_awready ;
wire  [DWID-1:0] slv12_wdata ;
wire  [WSTRB-1:0] slv12_wstrb ;
wire  slv12_wlast ;
wire  slv12_wvalid ;
reg  slv12_wready ;
reg  [IDWID-1:0] slv12_bid ;
reg  [1:0] slv12_bresp ;
reg  slv12_bvalid ;
wire  slv12_bready ;

initial slv12_arready = 0;
initial slv12_awready = 0;
initial slv12_rvalid = 0;
initial slv12_bvalid = 0;

reg  [2:0] slv13_awsize ; initial slv13_awsize = 0;
reg  [2:0] slv13_arsize ; initial slv13_arsize = 0;

wire  [IDWID-1:0] slv13_arid ;
wire  [31:0] slv13_araddr ;
wire  [7:0] slv13_arlen ;
wire  [EXTRAS-1:0] slv13_arextras ;
wire  [1:0] slv13_arburst ;
wire  slv13_arvalid ;
reg  slv13_arready ;
reg  [IDWID-1:0] slv13_rid ;
reg  [DWID-1:0] slv13_rdata ;
reg  [1:0] slv13_rresp ;
reg  slv13_rlast ;
reg  slv13_rvalid ;
wire  slv13_rready ;

wire  [IDWID-1:0] slv13_awid ;
wire  [31:0] slv13_awaddr ;
wire  [7:0] slv13_awlen ;
wire  [EXTRAS-1:0] slv13_awextras ;
wire  [1:0] slv13_awburst ;
wire  slv13_awvalid ;
reg  slv13_awready ;
wire  [DWID-1:0] slv13_wdata ;
wire  [WSTRB-1:0] slv13_wstrb ;
wire  slv13_wlast ;
wire  slv13_wvalid ;
reg  slv13_wready ;
reg  [IDWID-1:0] slv13_bid ;
reg  [1:0] slv13_bresp ;
reg  slv13_bvalid ;
wire  slv13_bready ;

initial slv13_arready = 0;
initial slv13_awready = 0;
initial slv13_rvalid = 0;
initial slv13_bvalid = 0;

reg  [2:0] slv14_awsize ; initial slv14_awsize = 0;
reg  [2:0] slv14_arsize ; initial slv14_arsize = 0;

wire  [IDWID-1:0] slv14_arid ;
wire  [31:0] slv14_araddr ;
wire  [7:0] slv14_arlen ;
wire  [EXTRAS-1:0] slv14_arextras ;
wire  [1:0] slv14_arburst ;
wire  slv14_arvalid ;
reg  slv14_arready ;
reg  [IDWID-1:0] slv14_rid ;
reg  [DWID-1:0] slv14_rdata ;
reg  [1:0] slv14_rresp ;
reg  slv14_rlast ;
reg  slv14_rvalid ;
wire  slv14_rready ;

wire  [IDWID-1:0] slv14_awid ;
wire  [31:0] slv14_awaddr ;
wire  [7:0] slv14_awlen ;
wire  [EXTRAS-1:0] slv14_awextras ;
wire  [1:0] slv14_awburst ;
wire  slv14_awvalid ;
reg  slv14_awready ;
wire  [DWID-1:0] slv14_wdata ;
wire  [WSTRB-1:0] slv14_wstrb ;
wire  slv14_wlast ;
wire  slv14_wvalid ;
reg  slv14_wready ;
reg  [IDWID-1:0] slv14_bid ;
reg  [1:0] slv14_bresp ;
reg  slv14_bvalid ;
wire  slv14_bready ;

initial slv14_arready = 0;
initial slv14_awready = 0;
initial slv14_rvalid = 0;
initial slv14_bvalid = 0;

reg  [2:0] slv15_awsize ; initial slv15_awsize = 0;
reg  [2:0] slv15_arsize ; initial slv15_arsize = 0;

wire  [IDWID-1:0] slv15_arid ;
wire  [31:0] slv15_araddr ;
wire  [7:0] slv15_arlen ;
wire  [EXTRAS-1:0] slv15_arextras ;
wire  [1:0] slv15_arburst ;
wire  slv15_arvalid ;
reg  slv15_arready ;
reg  [IDWID-1:0] slv15_rid ;
reg  [DWID-1:0] slv15_rdata ;
reg  [1:0] slv15_rresp ;
reg  slv15_rlast ;
reg  slv15_rvalid ;
wire  slv15_rready ;

wire  [IDWID-1:0] slv15_awid ;
wire  [31:0] slv15_awaddr ;
wire  [7:0] slv15_awlen ;
wire  [EXTRAS-1:0] slv15_awextras ;
wire  [1:0] slv15_awburst ;
wire  slv15_awvalid ;
reg  slv15_awready ;
wire  [DWID-1:0] slv15_wdata ;
wire  [WSTRB-1:0] slv15_wstrb ;
wire  slv15_wlast ;
wire  slv15_wvalid ;
reg  slv15_wready ;
reg  [IDWID-1:0] slv15_bid ;
reg  [1:0] slv15_bresp ;
reg  slv15_bvalid ;
wire  slv15_bready ;

initial slv15_arready = 0;
initial slv15_awready = 0;
initial slv15_rvalid = 0;
initial slv15_bvalid = 0;

reg  [2:0] slv2_awsize ; initial slv2_awsize = 0;
reg  [2:0] slv2_arsize ; initial slv2_arsize = 0;

wire  [IDWID-1:0] slv2_arid ;
wire  [31:0] slv2_araddr ;
wire  [7:0] slv2_arlen ;
wire  [EXTRAS-1:0] slv2_arextras ;
wire  [1:0] slv2_arburst ;
wire  slv2_arvalid ;
reg  slv2_arready ;
reg  [IDWID-1:0] slv2_rid ;
reg  [DWID-1:0] slv2_rdata ;
reg  [1:0] slv2_rresp ;
reg  slv2_rlast ;
reg  slv2_rvalid ;
wire  slv2_rready ;

wire  [IDWID-1:0] slv2_awid ;
wire  [31:0] slv2_awaddr ;
wire  [7:0] slv2_awlen ;
wire  [EXTRAS-1:0] slv2_awextras ;
wire  [1:0] slv2_awburst ;
wire  slv2_awvalid ;
reg  slv2_awready ;
wire  [DWID-1:0] slv2_wdata ;
wire  [WSTRB-1:0] slv2_wstrb ;
wire  slv2_wlast ;
wire  slv2_wvalid ;
reg  slv2_wready ;
reg  [IDWID-1:0] slv2_bid ;
reg  [1:0] slv2_bresp ;
reg  slv2_bvalid ;
wire  slv2_bready ;

initial slv2_arready = 0;
initial slv2_awready = 0;
initial slv2_rvalid = 0;
initial slv2_bvalid = 0;

reg  [2:0] slv3_awsize ; initial slv3_awsize = 0;
reg  [2:0] slv3_arsize ; initial slv3_arsize = 0;

wire  [IDWID-1:0] slv3_arid ;
wire  [31:0] slv3_araddr ;
wire  [7:0] slv3_arlen ;
wire  [EXTRAS-1:0] slv3_arextras ;
wire  [1:0] slv3_arburst ;
wire  slv3_arvalid ;
reg  slv3_arready ;
reg  [IDWID-1:0] slv3_rid ;
reg  [DWID-1:0] slv3_rdata ;
reg  [1:0] slv3_rresp ;
reg  slv3_rlast ;
reg  slv3_rvalid ;
wire  slv3_rready ;

wire  [IDWID-1:0] slv3_awid ;
wire  [31:0] slv3_awaddr ;
wire  [7:0] slv3_awlen ;
wire  [EXTRAS-1:0] slv3_awextras ;
wire  [1:0] slv3_awburst ;
wire  slv3_awvalid ;
reg  slv3_awready ;
wire  [DWID-1:0] slv3_wdata ;
wire  [WSTRB-1:0] slv3_wstrb ;
wire  slv3_wlast ;
wire  slv3_wvalid ;
reg  slv3_wready ;
reg  [IDWID-1:0] slv3_bid ;
reg  [1:0] slv3_bresp ;
reg  slv3_bvalid ;
wire  slv3_bready ;

initial slv3_arready = 0;
initial slv3_awready = 0;
initial slv3_rvalid = 0;
initial slv3_bvalid = 0;

reg  [2:0] slv4_awsize ; initial slv4_awsize = 0;
reg  [2:0] slv4_arsize ; initial slv4_arsize = 0;

wire  [IDWID-1:0] slv4_arid ;
wire  [31:0] slv4_araddr ;
wire  [7:0] slv4_arlen ;
wire  [EXTRAS-1:0] slv4_arextras ;
wire  [1:0] slv4_arburst ;
wire  slv4_arvalid ;
reg  slv4_arready ;
reg  [IDWID-1:0] slv4_rid ;
reg  [DWID-1:0] slv4_rdata ;
reg  [1:0] slv4_rresp ;
reg  slv4_rlast ;
reg  slv4_rvalid ;
wire  slv4_rready ;

wire  [IDWID-1:0] slv4_awid ;
wire  [31:0] slv4_awaddr ;
wire  [7:0] slv4_awlen ;
wire  [EXTRAS-1:0] slv4_awextras ;
wire  [1:0] slv4_awburst ;
wire  slv4_awvalid ;
reg  slv4_awready ;
wire  [DWID-1:0] slv4_wdata ;
wire  [WSTRB-1:0] slv4_wstrb ;
wire  slv4_wlast ;
wire  slv4_wvalid ;
reg  slv4_wready ;
reg  [IDWID-1:0] slv4_bid ;
reg  [1:0] slv4_bresp ;
reg  slv4_bvalid ;
wire  slv4_bready ;

initial slv4_arready = 0;
initial slv4_awready = 0;
initial slv4_rvalid = 0;
initial slv4_bvalid = 0;

reg  [2:0] slv5_awsize ; initial slv5_awsize = 0;
reg  [2:0] slv5_arsize ; initial slv5_arsize = 0;

wire  [IDWID-1:0] slv5_arid ;
wire  [31:0] slv5_araddr ;
wire  [7:0] slv5_arlen ;
wire  [EXTRAS-1:0] slv5_arextras ;
wire  [1:0] slv5_arburst ;
wire  slv5_arvalid ;
reg  slv5_arready ;
reg  [IDWID-1:0] slv5_rid ;
reg  [DWID-1:0] slv5_rdata ;
reg  [1:0] slv5_rresp ;
reg  slv5_rlast ;
reg  slv5_rvalid ;
wire  slv5_rready ;

wire  [IDWID-1:0] slv5_awid ;
wire  [31:0] slv5_awaddr ;
wire  [7:0] slv5_awlen ;
wire  [EXTRAS-1:0] slv5_awextras ;
wire  [1:0] slv5_awburst ;
wire  slv5_awvalid ;
reg  slv5_awready ;
wire  [DWID-1:0] slv5_wdata ;
wire  [WSTRB-1:0] slv5_wstrb ;
wire  slv5_wlast ;
wire  slv5_wvalid ;
reg  slv5_wready ;
reg  [IDWID-1:0] slv5_bid ;
reg  [1:0] slv5_bresp ;
reg  slv5_bvalid ;
wire  slv5_bready ;

initial slv5_arready = 0;
initial slv5_awready = 0;
initial slv5_rvalid = 0;
initial slv5_bvalid = 0;

reg  [2:0] slv6_awsize ; initial slv6_awsize = 0;
reg  [2:0] slv6_arsize ; initial slv6_arsize = 0;

wire  [IDWID-1:0] slv6_arid ;
wire  [31:0] slv6_araddr ;
wire  [7:0] slv6_arlen ;
wire  [EXTRAS-1:0] slv6_arextras ;
wire  [1:0] slv6_arburst ;
wire  slv6_arvalid ;
reg  slv6_arready ;
reg  [IDWID-1:0] slv6_rid ;
reg  [DWID-1:0] slv6_rdata ;
reg  [1:0] slv6_rresp ;
reg  slv6_rlast ;
reg  slv6_rvalid ;
wire  slv6_rready ;

wire  [IDWID-1:0] slv6_awid ;
wire  [31:0] slv6_awaddr ;
wire  [7:0] slv6_awlen ;
wire  [EXTRAS-1:0] slv6_awextras ;
wire  [1:0] slv6_awburst ;
wire  slv6_awvalid ;
reg  slv6_awready ;
wire  [DWID-1:0] slv6_wdata ;
wire  [WSTRB-1:0] slv6_wstrb ;
wire  slv6_wlast ;
wire  slv6_wvalid ;
reg  slv6_wready ;
reg  [IDWID-1:0] slv6_bid ;
reg  [1:0] slv6_bresp ;
reg  slv6_bvalid ;
wire  slv6_bready ;

initial slv6_arready = 0;
initial slv6_awready = 0;
initial slv6_rvalid = 0;
initial slv6_bvalid = 0;

reg  [2:0] slv7_awsize ; initial slv7_awsize = 0;
reg  [2:0] slv7_arsize ; initial slv7_arsize = 0;

wire  [IDWID-1:0] slv7_arid ;
wire  [31:0] slv7_araddr ;
wire  [7:0] slv7_arlen ;
wire  [EXTRAS-1:0] slv7_arextras ;
wire  [1:0] slv7_arburst ;
wire  slv7_arvalid ;
reg  slv7_arready ;
reg  [IDWID-1:0] slv7_rid ;
reg  [DWID-1:0] slv7_rdata ;
reg  [1:0] slv7_rresp ;
reg  slv7_rlast ;
reg  slv7_rvalid ;
wire  slv7_rready ;

wire  [IDWID-1:0] slv7_awid ;
wire  [31:0] slv7_awaddr ;
wire  [7:0] slv7_awlen ;
wire  [EXTRAS-1:0] slv7_awextras ;
wire  [1:0] slv7_awburst ;
wire  slv7_awvalid ;
reg  slv7_awready ;
wire  [DWID-1:0] slv7_wdata ;
wire  [WSTRB-1:0] slv7_wstrb ;
wire  slv7_wlast ;
wire  slv7_wvalid ;
reg  slv7_wready ;
reg  [IDWID-1:0] slv7_bid ;
reg  [1:0] slv7_bresp ;
reg  slv7_bvalid ;
wire  slv7_bready ;

initial slv7_arready = 0;
initial slv7_awready = 0;
initial slv7_rvalid = 0;
initial slv7_bvalid = 0;

reg  [2:0] slv8_awsize ; initial slv8_awsize = 0;
reg  [2:0] slv8_arsize ; initial slv8_arsize = 0;

wire  [IDWID-1:0] slv8_arid ;
wire  [31:0] slv8_araddr ;
wire  [7:0] slv8_arlen ;
wire  [EXTRAS-1:0] slv8_arextras ;
wire  [1:0] slv8_arburst ;
wire  slv8_arvalid ;
reg  slv8_arready ;
reg  [IDWID-1:0] slv8_rid ;
reg  [DWID-1:0] slv8_rdata ;
reg  [1:0] slv8_rresp ;
reg  slv8_rlast ;
reg  slv8_rvalid ;
wire  slv8_rready ;

wire  [IDWID-1:0] slv8_awid ;
wire  [31:0] slv8_awaddr ;
wire  [7:0] slv8_awlen ;
wire  [EXTRAS-1:0] slv8_awextras ;
wire  [1:0] slv8_awburst ;
wire  slv8_awvalid ;
reg  slv8_awready ;
wire  [DWID-1:0] slv8_wdata ;
wire  [WSTRB-1:0] slv8_wstrb ;
wire  slv8_wlast ;
wire  slv8_wvalid ;
reg  slv8_wready ;
reg  [IDWID-1:0] slv8_bid ;
reg  [1:0] slv8_bresp ;
reg  slv8_bvalid ;
wire  slv8_bready ;

initial slv8_arready = 0;
initial slv8_awready = 0;
initial slv8_rvalid = 0;
initial slv8_bvalid = 0;

reg  [2:0] slv9_awsize ; initial slv9_awsize = 0;
reg  [2:0] slv9_arsize ; initial slv9_arsize = 0;

wire  [IDWID-1:0] slv9_arid ;
wire  [31:0] slv9_araddr ;
wire  [7:0] slv9_arlen ;
wire  [EXTRAS-1:0] slv9_arextras ;
wire  [1:0] slv9_arburst ;
wire  slv9_arvalid ;
reg  slv9_arready ;
reg  [IDWID-1:0] slv9_rid ;
reg  [DWID-1:0] slv9_rdata ;
reg  [1:0] slv9_rresp ;
reg  slv9_rlast ;
reg  slv9_rvalid ;
wire  slv9_rready ;

wire  [IDWID-1:0] slv9_awid ;
wire  [31:0] slv9_awaddr ;
wire  [7:0] slv9_awlen ;
wire  [EXTRAS-1:0] slv9_awextras ;
wire  [1:0] slv9_awburst ;
wire  slv9_awvalid ;
reg  slv9_awready ;
wire  [DWID-1:0] slv9_wdata ;
wire  [WSTRB-1:0] slv9_wstrb ;
wire  slv9_wlast ;
wire  slv9_wvalid ;
reg  slv9_wready ;
reg  [IDWID-1:0] slv9_bid ;
reg  [1:0] slv9_bresp ;
reg  slv9_bvalid ;
wire  slv9_bready ;

initial slv9_arready = 0;
initial slv9_awready = 0;
initial slv9_rvalid = 0;
initial slv9_bvalid = 0;

reg  [2:0] mst0_awsize ; initial mst0_awsize = 0;
reg  [2:0] mst0_arsize ; initial mst0_arsize = 0;

reg  [IDWID-1:0] mst0_arid ;
reg  [31:0] mst0_araddr ;
reg  [7:0] mst0_arlen ;
reg  [EXTRAS-1:0] mst0_arextras ;
reg  [1:0] mst0_arburst ;
reg  mst0_arvalid ;
wire  mst0_arready ;
wire  [IDWID-1:0] mst0_rid ;
wire  [DWID-1:0] mst0_rdata ;
wire  [1:0] mst0_rresp ;
wire  mst0_rlast ;
wire  mst0_rvalid ;
reg  mst0_rready ;

reg  [IDWID-1:0] mst0_awid ;
reg  [31:0] mst0_awaddr ;
reg  [7:0] mst0_awlen ;
reg  [EXTRAS-1:0] mst0_awextras ;
reg  [1:0] mst0_awburst ;
reg  mst0_awvalid ;
wire  mst0_awready ;
reg  [DWID-1:0] mst0_wdata ;
reg  [WSTRB-1:0] mst0_wstrb ;
reg  mst0_wlast ;
reg  mst0_wvalid ;
wire  mst0_wready ;
wire  [IDWID-1:0] mst0_bid ;
wire  [1:0] mst0_bresp ;
wire  mst0_bvalid ;
reg  mst0_bready ;

initial mst0_bready = 0;
initial mst0_wvalid = 0;
initial mst0_arvalid = 0;
initial mst0_awvalid = 0;
initial mst0_rready = 0;

reg  [2:0] mst1_awsize ; initial mst1_awsize = 0;
reg  [2:0] mst1_arsize ; initial mst1_arsize = 0;

reg  [IDWID-1:0] mst1_arid ;
reg  [31:0] mst1_araddr ;
reg  [7:0] mst1_arlen ;
reg  [EXTRAS-1:0] mst1_arextras ;
reg  [1:0] mst1_arburst ;
reg  mst1_arvalid ;
wire  mst1_arready ;
wire  [IDWID-1:0] mst1_rid ;
wire  [DWID-1:0] mst1_rdata ;
wire  [1:0] mst1_rresp ;
wire  mst1_rlast ;
wire  mst1_rvalid ;
reg  mst1_rready ;

reg  [IDWID-1:0] mst1_awid ;
reg  [31:0] mst1_awaddr ;
reg  [7:0] mst1_awlen ;
reg  [EXTRAS-1:0] mst1_awextras ;
reg  [1:0] mst1_awburst ;
reg  mst1_awvalid ;
wire  mst1_awready ;
reg  [DWID-1:0] mst1_wdata ;
reg  [WSTRB-1:0] mst1_wstrb ;
reg  mst1_wlast ;
reg  mst1_wvalid ;
wire  mst1_wready ;
wire  [IDWID-1:0] mst1_bid ;
wire  [1:0] mst1_bresp ;
wire  mst1_bvalid ;
reg  mst1_bready ;

initial mst1_bready = 0;
initial mst1_wvalid = 0;
initial mst1_arvalid = 0;
initial mst1_awvalid = 0;
initial mst1_rready = 0;

reg  [2:0] mst10_awsize ; initial mst10_awsize = 0;
reg  [2:0] mst10_arsize ; initial mst10_arsize = 0;

reg  [IDWID-1:0] mst10_arid ;
reg  [31:0] mst10_araddr ;
reg  [7:0] mst10_arlen ;
reg  [EXTRAS-1:0] mst10_arextras ;
reg  [1:0] mst10_arburst ;
reg  mst10_arvalid ;
wire  mst10_arready ;
wire  [IDWID-1:0] mst10_rid ;
wire  [DWID-1:0] mst10_rdata ;
wire  [1:0] mst10_rresp ;
wire  mst10_rlast ;
wire  mst10_rvalid ;
reg  mst10_rready ;

reg  [IDWID-1:0] mst10_awid ;
reg  [31:0] mst10_awaddr ;
reg  [7:0] mst10_awlen ;
reg  [EXTRAS-1:0] mst10_awextras ;
reg  [1:0] mst10_awburst ;
reg  mst10_awvalid ;
wire  mst10_awready ;
reg  [DWID-1:0] mst10_wdata ;
reg  [WSTRB-1:0] mst10_wstrb ;
reg  mst10_wlast ;
reg  mst10_wvalid ;
wire  mst10_wready ;
wire  [IDWID-1:0] mst10_bid ;
wire  [1:0] mst10_bresp ;
wire  mst10_bvalid ;
reg  mst10_bready ;

initial mst10_bready = 0;
initial mst10_wvalid = 0;
initial mst10_arvalid = 0;
initial mst10_awvalid = 0;
initial mst10_rready = 0;

reg  [2:0] mst11_awsize ; initial mst11_awsize = 0;
reg  [2:0] mst11_arsize ; initial mst11_arsize = 0;

reg  [IDWID-1:0] mst11_arid ;
reg  [31:0] mst11_araddr ;
reg  [7:0] mst11_arlen ;
reg  [EXTRAS-1:0] mst11_arextras ;
reg  [1:0] mst11_arburst ;
reg  mst11_arvalid ;
wire  mst11_arready ;
wire  [IDWID-1:0] mst11_rid ;
wire  [DWID-1:0] mst11_rdata ;
wire  [1:0] mst11_rresp ;
wire  mst11_rlast ;
wire  mst11_rvalid ;
reg  mst11_rready ;

reg  [IDWID-1:0] mst11_awid ;
reg  [31:0] mst11_awaddr ;
reg  [7:0] mst11_awlen ;
reg  [EXTRAS-1:0] mst11_awextras ;
reg  [1:0] mst11_awburst ;
reg  mst11_awvalid ;
wire  mst11_awready ;
reg  [DWID-1:0] mst11_wdata ;
reg  [WSTRB-1:0] mst11_wstrb ;
reg  mst11_wlast ;
reg  mst11_wvalid ;
wire  mst11_wready ;
wire  [IDWID-1:0] mst11_bid ;
wire  [1:0] mst11_bresp ;
wire  mst11_bvalid ;
reg  mst11_bready ;

initial mst11_bready = 0;
initial mst11_wvalid = 0;
initial mst11_arvalid = 0;
initial mst11_awvalid = 0;
initial mst11_rready = 0;

reg  [2:0] mst12_awsize ; initial mst12_awsize = 0;
reg  [2:0] mst12_arsize ; initial mst12_arsize = 0;

reg  [IDWID-1:0] mst12_arid ;
reg  [31:0] mst12_araddr ;
reg  [7:0] mst12_arlen ;
reg  [EXTRAS-1:0] mst12_arextras ;
reg  [1:0] mst12_arburst ;
reg  mst12_arvalid ;
wire  mst12_arready ;
wire  [IDWID-1:0] mst12_rid ;
wire  [DWID-1:0] mst12_rdata ;
wire  [1:0] mst12_rresp ;
wire  mst12_rlast ;
wire  mst12_rvalid ;
reg  mst12_rready ;

reg  [IDWID-1:0] mst12_awid ;
reg  [31:0] mst12_awaddr ;
reg  [7:0] mst12_awlen ;
reg  [EXTRAS-1:0] mst12_awextras ;
reg  [1:0] mst12_awburst ;
reg  mst12_awvalid ;
wire  mst12_awready ;
reg  [DWID-1:0] mst12_wdata ;
reg  [WSTRB-1:0] mst12_wstrb ;
reg  mst12_wlast ;
reg  mst12_wvalid ;
wire  mst12_wready ;
wire  [IDWID-1:0] mst12_bid ;
wire  [1:0] mst12_bresp ;
wire  mst12_bvalid ;
reg  mst12_bready ;

initial mst12_bready = 0;
initial mst12_wvalid = 0;
initial mst12_arvalid = 0;
initial mst12_awvalid = 0;
initial mst12_rready = 0;

reg  [2:0] mst13_awsize ; initial mst13_awsize = 0;
reg  [2:0] mst13_arsize ; initial mst13_arsize = 0;

reg  [IDWID-1:0] mst13_arid ;
reg  [31:0] mst13_araddr ;
reg  [7:0] mst13_arlen ;
reg  [EXTRAS-1:0] mst13_arextras ;
reg  [1:0] mst13_arburst ;
reg  mst13_arvalid ;
wire  mst13_arready ;
wire  [IDWID-1:0] mst13_rid ;
wire  [DWID-1:0] mst13_rdata ;
wire  [1:0] mst13_rresp ;
wire  mst13_rlast ;
wire  mst13_rvalid ;
reg  mst13_rready ;

reg  [IDWID-1:0] mst13_awid ;
reg  [31:0] mst13_awaddr ;
reg  [7:0] mst13_awlen ;
reg  [EXTRAS-1:0] mst13_awextras ;
reg  [1:0] mst13_awburst ;
reg  mst13_awvalid ;
wire  mst13_awready ;
reg  [DWID-1:0] mst13_wdata ;
reg  [WSTRB-1:0] mst13_wstrb ;
reg  mst13_wlast ;
reg  mst13_wvalid ;
wire  mst13_wready ;
wire  [IDWID-1:0] mst13_bid ;
wire  [1:0] mst13_bresp ;
wire  mst13_bvalid ;
reg  mst13_bready ;

initial mst13_bready = 0;
initial mst13_wvalid = 0;
initial mst13_arvalid = 0;
initial mst13_awvalid = 0;
initial mst13_rready = 0;

reg  [2:0] mst14_awsize ; initial mst14_awsize = 0;
reg  [2:0] mst14_arsize ; initial mst14_arsize = 0;

reg  [IDWID-1:0] mst14_arid ;
reg  [31:0] mst14_araddr ;
reg  [7:0] mst14_arlen ;
reg  [EXTRAS-1:0] mst14_arextras ;
reg  [1:0] mst14_arburst ;
reg  mst14_arvalid ;
wire  mst14_arready ;
wire  [IDWID-1:0] mst14_rid ;
wire  [DWID-1:0] mst14_rdata ;
wire  [1:0] mst14_rresp ;
wire  mst14_rlast ;
wire  mst14_rvalid ;
reg  mst14_rready ;

reg  [IDWID-1:0] mst14_awid ;
reg  [31:0] mst14_awaddr ;
reg  [7:0] mst14_awlen ;
reg  [EXTRAS-1:0] mst14_awextras ;
reg  [1:0] mst14_awburst ;
reg  mst14_awvalid ;
wire  mst14_awready ;
reg  [DWID-1:0] mst14_wdata ;
reg  [WSTRB-1:0] mst14_wstrb ;
reg  mst14_wlast ;
reg  mst14_wvalid ;
wire  mst14_wready ;
wire  [IDWID-1:0] mst14_bid ;
wire  [1:0] mst14_bresp ;
wire  mst14_bvalid ;
reg  mst14_bready ;

initial mst14_bready = 0;
initial mst14_wvalid = 0;
initial mst14_arvalid = 0;
initial mst14_awvalid = 0;
initial mst14_rready = 0;

reg  [2:0] mst15_awsize ; initial mst15_awsize = 0;
reg  [2:0] mst15_arsize ; initial mst15_arsize = 0;

reg  [IDWID-1:0] mst15_arid ;
reg  [31:0] mst15_araddr ;
reg  [7:0] mst15_arlen ;
reg  [EXTRAS-1:0] mst15_arextras ;
reg  [1:0] mst15_arburst ;
reg  mst15_arvalid ;
wire  mst15_arready ;
wire  [IDWID-1:0] mst15_rid ;
wire  [DWID-1:0] mst15_rdata ;
wire  [1:0] mst15_rresp ;
wire  mst15_rlast ;
wire  mst15_rvalid ;
reg  mst15_rready ;

reg  [IDWID-1:0] mst15_awid ;
reg  [31:0] mst15_awaddr ;
reg  [7:0] mst15_awlen ;
reg  [EXTRAS-1:0] mst15_awextras ;
reg  [1:0] mst15_awburst ;
reg  mst15_awvalid ;
wire  mst15_awready ;
reg  [DWID-1:0] mst15_wdata ;
reg  [WSTRB-1:0] mst15_wstrb ;
reg  mst15_wlast ;
reg  mst15_wvalid ;
wire  mst15_wready ;
wire  [IDWID-1:0] mst15_bid ;
wire  [1:0] mst15_bresp ;
wire  mst15_bvalid ;
reg  mst15_bready ;

initial mst15_bready = 0;
initial mst15_wvalid = 0;
initial mst15_arvalid = 0;
initial mst15_awvalid = 0;
initial mst15_rready = 0;

reg  [2:0] mst2_awsize ; initial mst2_awsize = 0;
reg  [2:0] mst2_arsize ; initial mst2_arsize = 0;

reg  [IDWID-1:0] mst2_arid ;
reg  [31:0] mst2_araddr ;
reg  [7:0] mst2_arlen ;
reg  [EXTRAS-1:0] mst2_arextras ;
reg  [1:0] mst2_arburst ;
reg  mst2_arvalid ;
wire  mst2_arready ;
wire  [IDWID-1:0] mst2_rid ;
wire  [DWID-1:0] mst2_rdata ;
wire  [1:0] mst2_rresp ;
wire  mst2_rlast ;
wire  mst2_rvalid ;
reg  mst2_rready ;

reg  [IDWID-1:0] mst2_awid ;
reg  [31:0] mst2_awaddr ;
reg  [7:0] mst2_awlen ;
reg  [EXTRAS-1:0] mst2_awextras ;
reg  [1:0] mst2_awburst ;
reg  mst2_awvalid ;
wire  mst2_awready ;
reg  [DWID-1:0] mst2_wdata ;
reg  [WSTRB-1:0] mst2_wstrb ;
reg  mst2_wlast ;
reg  mst2_wvalid ;
wire  mst2_wready ;
wire  [IDWID-1:0] mst2_bid ;
wire  [1:0] mst2_bresp ;
wire  mst2_bvalid ;
reg  mst2_bready ;

initial mst2_bready = 0;
initial mst2_wvalid = 0;
initial mst2_arvalid = 0;
initial mst2_awvalid = 0;
initial mst2_rready = 0;

reg  [2:0] mst3_awsize ; initial mst3_awsize = 0;
reg  [2:0] mst3_arsize ; initial mst3_arsize = 0;

reg  [IDWID-1:0] mst3_arid ;
reg  [31:0] mst3_araddr ;
reg  [7:0] mst3_arlen ;
reg  [EXTRAS-1:0] mst3_arextras ;
reg  [1:0] mst3_arburst ;
reg  mst3_arvalid ;
wire  mst3_arready ;
wire  [IDWID-1:0] mst3_rid ;
wire  [DWID-1:0] mst3_rdata ;
wire  [1:0] mst3_rresp ;
wire  mst3_rlast ;
wire  mst3_rvalid ;
reg  mst3_rready ;

reg  [IDWID-1:0] mst3_awid ;
reg  [31:0] mst3_awaddr ;
reg  [7:0] mst3_awlen ;
reg  [EXTRAS-1:0] mst3_awextras ;
reg  [1:0] mst3_awburst ;
reg  mst3_awvalid ;
wire  mst3_awready ;
reg  [DWID-1:0] mst3_wdata ;
reg  [WSTRB-1:0] mst3_wstrb ;
reg  mst3_wlast ;
reg  mst3_wvalid ;
wire  mst3_wready ;
wire  [IDWID-1:0] mst3_bid ;
wire  [1:0] mst3_bresp ;
wire  mst3_bvalid ;
reg  mst3_bready ;

initial mst3_bready = 0;
initial mst3_wvalid = 0;
initial mst3_arvalid = 0;
initial mst3_awvalid = 0;
initial mst3_rready = 0;

reg  [2:0] mst4_awsize ; initial mst4_awsize = 0;
reg  [2:0] mst4_arsize ; initial mst4_arsize = 0;

reg  [IDWID-1:0] mst4_arid ;
reg  [31:0] mst4_araddr ;
reg  [7:0] mst4_arlen ;
reg  [EXTRAS-1:0] mst4_arextras ;
reg  [1:0] mst4_arburst ;
reg  mst4_arvalid ;
wire  mst4_arready ;
wire  [IDWID-1:0] mst4_rid ;
wire  [DWID-1:0] mst4_rdata ;
wire  [1:0] mst4_rresp ;
wire  mst4_rlast ;
wire  mst4_rvalid ;
reg  mst4_rready ;

reg  [IDWID-1:0] mst4_awid ;
reg  [31:0] mst4_awaddr ;
reg  [7:0] mst4_awlen ;
reg  [EXTRAS-1:0] mst4_awextras ;
reg  [1:0] mst4_awburst ;
reg  mst4_awvalid ;
wire  mst4_awready ;
reg  [DWID-1:0] mst4_wdata ;
reg  [WSTRB-1:0] mst4_wstrb ;
reg  mst4_wlast ;
reg  mst4_wvalid ;
wire  mst4_wready ;
wire  [IDWID-1:0] mst4_bid ;
wire  [1:0] mst4_bresp ;
wire  mst4_bvalid ;
reg  mst4_bready ;

initial mst4_bready = 0;
initial mst4_wvalid = 0;
initial mst4_arvalid = 0;
initial mst4_awvalid = 0;
initial mst4_rready = 0;

reg  [2:0] mst5_awsize ; initial mst5_awsize = 0;
reg  [2:0] mst5_arsize ; initial mst5_arsize = 0;

reg  [IDWID-1:0] mst5_arid ;
reg  [31:0] mst5_araddr ;
reg  [7:0] mst5_arlen ;
reg  [EXTRAS-1:0] mst5_arextras ;
reg  [1:0] mst5_arburst ;
reg  mst5_arvalid ;
wire  mst5_arready ;
wire  [IDWID-1:0] mst5_rid ;
wire  [DWID-1:0] mst5_rdata ;
wire  [1:0] mst5_rresp ;
wire  mst5_rlast ;
wire  mst5_rvalid ;
reg  mst5_rready ;

reg  [IDWID-1:0] mst5_awid ;
reg  [31:0] mst5_awaddr ;
reg  [7:0] mst5_awlen ;
reg  [EXTRAS-1:0] mst5_awextras ;
reg  [1:0] mst5_awburst ;
reg  mst5_awvalid ;
wire  mst5_awready ;
reg  [DWID-1:0] mst5_wdata ;
reg  [WSTRB-1:0] mst5_wstrb ;
reg  mst5_wlast ;
reg  mst5_wvalid ;
wire  mst5_wready ;
wire  [IDWID-1:0] mst5_bid ;
wire  [1:0] mst5_bresp ;
wire  mst5_bvalid ;
reg  mst5_bready ;

initial mst5_bready = 0;
initial mst5_wvalid = 0;
initial mst5_arvalid = 0;
initial mst5_awvalid = 0;
initial mst5_rready = 0;

reg  [2:0] mst6_awsize ; initial mst6_awsize = 0;
reg  [2:0] mst6_arsize ; initial mst6_arsize = 0;

reg  [IDWID-1:0] mst6_arid ;
reg  [31:0] mst6_araddr ;
reg  [7:0] mst6_arlen ;
reg  [EXTRAS-1:0] mst6_arextras ;
reg  [1:0] mst6_arburst ;
reg  mst6_arvalid ;
wire  mst6_arready ;
wire  [IDWID-1:0] mst6_rid ;
wire  [DWID-1:0] mst6_rdata ;
wire  [1:0] mst6_rresp ;
wire  mst6_rlast ;
wire  mst6_rvalid ;
reg  mst6_rready ;

reg  [IDWID-1:0] mst6_awid ;
reg  [31:0] mst6_awaddr ;
reg  [7:0] mst6_awlen ;
reg  [EXTRAS-1:0] mst6_awextras ;
reg  [1:0] mst6_awburst ;
reg  mst6_awvalid ;
wire  mst6_awready ;
reg  [DWID-1:0] mst6_wdata ;
reg  [WSTRB-1:0] mst6_wstrb ;
reg  mst6_wlast ;
reg  mst6_wvalid ;
wire  mst6_wready ;
wire  [IDWID-1:0] mst6_bid ;
wire  [1:0] mst6_bresp ;
wire  mst6_bvalid ;
reg  mst6_bready ;

initial mst6_bready = 0;
initial mst6_wvalid = 0;
initial mst6_arvalid = 0;
initial mst6_awvalid = 0;
initial mst6_rready = 0;

reg  [2:0] mst7_awsize ; initial mst7_awsize = 0;
reg  [2:0] mst7_arsize ; initial mst7_arsize = 0;

reg  [IDWID-1:0] mst7_arid ;
reg  [31:0] mst7_araddr ;
reg  [7:0] mst7_arlen ;
reg  [EXTRAS-1:0] mst7_arextras ;
reg  [1:0] mst7_arburst ;
reg  mst7_arvalid ;
wire  mst7_arready ;
wire  [IDWID-1:0] mst7_rid ;
wire  [DWID-1:0] mst7_rdata ;
wire  [1:0] mst7_rresp ;
wire  mst7_rlast ;
wire  mst7_rvalid ;
reg  mst7_rready ;

reg  [IDWID-1:0] mst7_awid ;
reg  [31:0] mst7_awaddr ;
reg  [7:0] mst7_awlen ;
reg  [EXTRAS-1:0] mst7_awextras ;
reg  [1:0] mst7_awburst ;
reg  mst7_awvalid ;
wire  mst7_awready ;
reg  [DWID-1:0] mst7_wdata ;
reg  [WSTRB-1:0] mst7_wstrb ;
reg  mst7_wlast ;
reg  mst7_wvalid ;
wire  mst7_wready ;
wire  [IDWID-1:0] mst7_bid ;
wire  [1:0] mst7_bresp ;
wire  mst7_bvalid ;
reg  mst7_bready ;

initial mst7_bready = 0;
initial mst7_wvalid = 0;
initial mst7_arvalid = 0;
initial mst7_awvalid = 0;
initial mst7_rready = 0;

reg  [2:0] mst8_awsize ; initial mst8_awsize = 0;
reg  [2:0] mst8_arsize ; initial mst8_arsize = 0;

reg  [IDWID-1:0] mst8_arid ;
reg  [31:0] mst8_araddr ;
reg  [7:0] mst8_arlen ;
reg  [EXTRAS-1:0] mst8_arextras ;
reg  [1:0] mst8_arburst ;
reg  mst8_arvalid ;
wire  mst8_arready ;
wire  [IDWID-1:0] mst8_rid ;
wire  [DWID-1:0] mst8_rdata ;
wire  [1:0] mst8_rresp ;
wire  mst8_rlast ;
wire  mst8_rvalid ;
reg  mst8_rready ;

reg  [IDWID-1:0] mst8_awid ;
reg  [31:0] mst8_awaddr ;
reg  [7:0] mst8_awlen ;
reg  [EXTRAS-1:0] mst8_awextras ;
reg  [1:0] mst8_awburst ;
reg  mst8_awvalid ;
wire  mst8_awready ;
reg  [DWID-1:0] mst8_wdata ;
reg  [WSTRB-1:0] mst8_wstrb ;
reg  mst8_wlast ;
reg  mst8_wvalid ;
wire  mst8_wready ;
wire  [IDWID-1:0] mst8_bid ;
wire  [1:0] mst8_bresp ;
wire  mst8_bvalid ;
reg  mst8_bready ;

initial mst8_bready = 0;
initial mst8_wvalid = 0;
initial mst8_arvalid = 0;
initial mst8_awvalid = 0;
initial mst8_rready = 0;

reg  [2:0] mst9_awsize ; initial mst9_awsize = 0;
reg  [2:0] mst9_arsize ; initial mst9_arsize = 0;

reg  [IDWID-1:0] mst9_arid ;
reg  [31:0] mst9_araddr ;
reg  [7:0] mst9_arlen ;
reg  [EXTRAS-1:0] mst9_arextras ;
reg  [1:0] mst9_arburst ;
reg  mst9_arvalid ;
wire  mst9_arready ;
wire  [IDWID-1:0] mst9_rid ;
wire  [DWID-1:0] mst9_rdata ;
wire  [1:0] mst9_rresp ;
wire  mst9_rlast ;
wire  mst9_rvalid ;
reg  mst9_rready ;

reg  [IDWID-1:0] mst9_awid ;
reg  [31:0] mst9_awaddr ;
reg  [7:0] mst9_awlen ;
reg  [EXTRAS-1:0] mst9_awextras ;
reg  [1:0] mst9_awburst ;
reg  mst9_awvalid ;
wire  mst9_awready ;
reg  [DWID-1:0] mst9_wdata ;
reg  [WSTRB-1:0] mst9_wstrb ;
reg  mst9_wlast ;
reg  mst9_wvalid ;
wire  mst9_wready ;
wire  [IDWID-1:0] mst9_bid ;
wire  [1:0] mst9_bresp ;
wire  mst9_bvalid ;
reg  mst9_bready ;

initial mst9_bready = 0;
initial mst9_wvalid = 0;
initial mst9_arvalid = 0;
initial mst9_awvalid = 0;
initial mst9_rready = 0;
x16 dut ( .clk(clk),.rst_n(rst_n)

    ,.slv0_araddr(slv0_araddr[31:0])
    ,.slv0_arburst(slv0_arburst[1:0])
    ,.slv0_arextras(slv0_arextras[(EXTRAS - 1):0])
    ,.slv0_arid(slv0_arid[(IDWID - 1):0])
    ,.slv0_arlen(slv0_arlen[7:0])
    ,.slv0_arready(slv0_arready)
    ,.slv0_arvalid(slv0_arvalid)
    ,.slv0_awaddr(slv0_awaddr[31:0])
    ,.slv0_awburst(slv0_awburst[1:0])
    ,.slv0_awextras(slv0_awextras[(EXTRAS - 1):0])
    ,.slv0_awid(slv0_awid[(IDWID - 1):0])
    ,.slv0_awlen(slv0_awlen[7:0])
    ,.slv0_awready(slv0_awready)
    ,.slv0_awvalid(slv0_awvalid)
    ,.slv0_bid(slv0_bid[(IDWID - 1):0])
    ,.slv0_bready(slv0_bready)
    ,.slv0_bresp(slv0_bresp[1:0])
    ,.slv0_bvalid(slv0_bvalid)
    ,.slv0_rdata(slv0_rdata[(DWID - 1):0])
    ,.slv0_rid(slv0_rid[(IDWID - 1):0])
    ,.slv0_rlast(slv0_rlast)
    ,.slv0_rready(slv0_rready)
    ,.slv0_rresp(slv0_rresp[1:0])
    ,.slv0_rvalid(slv0_rvalid)
    ,.slv0_wdata(slv0_wdata[(DWID - 1):0])
    ,.slv0_wlast(slv0_wlast)
    ,.slv0_wready(slv0_wready)
    ,.slv0_wstrb(slv0_wstrb[(WSTRB - 1):0])
    ,.slv0_wvalid(slv0_wvalid)


    ,.slv1_araddr(slv1_araddr[31:0])
    ,.slv1_arburst(slv1_arburst[1:0])
    ,.slv1_arextras(slv1_arextras[(EXTRAS - 1):0])
    ,.slv1_arid(slv1_arid[(IDWID - 1):0])
    ,.slv1_arlen(slv1_arlen[7:0])
    ,.slv1_arready(slv1_arready)
    ,.slv1_arvalid(slv1_arvalid)
    ,.slv1_awaddr(slv1_awaddr[31:0])
    ,.slv1_awburst(slv1_awburst[1:0])
    ,.slv1_awextras(slv1_awextras[(EXTRAS - 1):0])
    ,.slv1_awid(slv1_awid[(IDWID - 1):0])
    ,.slv1_awlen(slv1_awlen[7:0])
    ,.slv1_awready(slv1_awready)
    ,.slv1_awvalid(slv1_awvalid)
    ,.slv1_bid(slv1_bid[(IDWID - 1):0])
    ,.slv1_bready(slv1_bready)
    ,.slv1_bresp(slv1_bresp[1:0])
    ,.slv1_bvalid(slv1_bvalid)
    ,.slv1_rdata(slv1_rdata[(DWID - 1):0])
    ,.slv1_rid(slv1_rid[(IDWID - 1):0])
    ,.slv1_rlast(slv1_rlast)
    ,.slv1_rready(slv1_rready)
    ,.slv1_rresp(slv1_rresp[1:0])
    ,.slv1_rvalid(slv1_rvalid)
    ,.slv1_wdata(slv1_wdata[(DWID - 1):0])
    ,.slv1_wlast(slv1_wlast)
    ,.slv1_wready(slv1_wready)
    ,.slv1_wstrb(slv1_wstrb[(WSTRB - 1):0])
    ,.slv1_wvalid(slv1_wvalid)


    ,.slv10_araddr(slv10_araddr[31:0])
    ,.slv10_arburst(slv10_arburst[1:0])
    ,.slv10_arextras(slv10_arextras[(EXTRAS - 1):0])
    ,.slv10_arid(slv10_arid[(IDWID - 1):0])
    ,.slv10_arlen(slv10_arlen[7:0])
    ,.slv10_arready(slv10_arready)
    ,.slv10_arvalid(slv10_arvalid)
    ,.slv10_awaddr(slv10_awaddr[31:0])
    ,.slv10_awburst(slv10_awburst[1:0])
    ,.slv10_awextras(slv10_awextras[(EXTRAS - 1):0])
    ,.slv10_awid(slv10_awid[(IDWID - 1):0])
    ,.slv10_awlen(slv10_awlen[7:0])
    ,.slv10_awready(slv10_awready)
    ,.slv10_awvalid(slv10_awvalid)
    ,.slv10_bid(slv10_bid[(IDWID - 1):0])
    ,.slv10_bready(slv10_bready)
    ,.slv10_bresp(slv10_bresp[1:0])
    ,.slv10_bvalid(slv10_bvalid)
    ,.slv10_rdata(slv10_rdata[(DWID - 1):0])
    ,.slv10_rid(slv10_rid[(IDWID - 1):0])
    ,.slv10_rlast(slv10_rlast)
    ,.slv10_rready(slv10_rready)
    ,.slv10_rresp(slv10_rresp[1:0])
    ,.slv10_rvalid(slv10_rvalid)
    ,.slv10_wdata(slv10_wdata[(DWID - 1):0])
    ,.slv10_wlast(slv10_wlast)
    ,.slv10_wready(slv10_wready)
    ,.slv10_wstrb(slv10_wstrb[(WSTRB - 1):0])
    ,.slv10_wvalid(slv10_wvalid)


    ,.slv11_araddr(slv11_araddr[31:0])
    ,.slv11_arburst(slv11_arburst[1:0])
    ,.slv11_arextras(slv11_arextras[(EXTRAS - 1):0])
    ,.slv11_arid(slv11_arid[(IDWID - 1):0])
    ,.slv11_arlen(slv11_arlen[7:0])
    ,.slv11_arready(slv11_arready)
    ,.slv11_arvalid(slv11_arvalid)
    ,.slv11_awaddr(slv11_awaddr[31:0])
    ,.slv11_awburst(slv11_awburst[1:0])
    ,.slv11_awextras(slv11_awextras[(EXTRAS - 1):0])
    ,.slv11_awid(slv11_awid[(IDWID - 1):0])
    ,.slv11_awlen(slv11_awlen[7:0])
    ,.slv11_awready(slv11_awready)
    ,.slv11_awvalid(slv11_awvalid)
    ,.slv11_bid(slv11_bid[(IDWID - 1):0])
    ,.slv11_bready(slv11_bready)
    ,.slv11_bresp(slv11_bresp[1:0])
    ,.slv11_bvalid(slv11_bvalid)
    ,.slv11_rdata(slv11_rdata[(DWID - 1):0])
    ,.slv11_rid(slv11_rid[(IDWID - 1):0])
    ,.slv11_rlast(slv11_rlast)
    ,.slv11_rready(slv11_rready)
    ,.slv11_rresp(slv11_rresp[1:0])
    ,.slv11_rvalid(slv11_rvalid)
    ,.slv11_wdata(slv11_wdata[(DWID - 1):0])
    ,.slv11_wlast(slv11_wlast)
    ,.slv11_wready(slv11_wready)
    ,.slv11_wstrb(slv11_wstrb[(WSTRB - 1):0])
    ,.slv11_wvalid(slv11_wvalid)


    ,.slv12_araddr(slv12_araddr[31:0])
    ,.slv12_arburst(slv12_arburst[1:0])
    ,.slv12_arextras(slv12_arextras[(EXTRAS - 1):0])
    ,.slv12_arid(slv12_arid[(IDWID - 1):0])
    ,.slv12_arlen(slv12_arlen[7:0])
    ,.slv12_arready(slv12_arready)
    ,.slv12_arvalid(slv12_arvalid)
    ,.slv12_awaddr(slv12_awaddr[31:0])
    ,.slv12_awburst(slv12_awburst[1:0])
    ,.slv12_awextras(slv12_awextras[(EXTRAS - 1):0])
    ,.slv12_awid(slv12_awid[(IDWID - 1):0])
    ,.slv12_awlen(slv12_awlen[7:0])
    ,.slv12_awready(slv12_awready)
    ,.slv12_awvalid(slv12_awvalid)
    ,.slv12_bid(slv12_bid[(IDWID - 1):0])
    ,.slv12_bready(slv12_bready)
    ,.slv12_bresp(slv12_bresp[1:0])
    ,.slv12_bvalid(slv12_bvalid)
    ,.slv12_rdata(slv12_rdata[(DWID - 1):0])
    ,.slv12_rid(slv12_rid[(IDWID - 1):0])
    ,.slv12_rlast(slv12_rlast)
    ,.slv12_rready(slv12_rready)
    ,.slv12_rresp(slv12_rresp[1:0])
    ,.slv12_rvalid(slv12_rvalid)
    ,.slv12_wdata(slv12_wdata[(DWID - 1):0])
    ,.slv12_wlast(slv12_wlast)
    ,.slv12_wready(slv12_wready)
    ,.slv12_wstrb(slv12_wstrb[(WSTRB - 1):0])
    ,.slv12_wvalid(slv12_wvalid)


    ,.slv13_araddr(slv13_araddr[31:0])
    ,.slv13_arburst(slv13_arburst[1:0])
    ,.slv13_arextras(slv13_arextras[(EXTRAS - 1):0])
    ,.slv13_arid(slv13_arid[(IDWID - 1):0])
    ,.slv13_arlen(slv13_arlen[7:0])
    ,.slv13_arready(slv13_arready)
    ,.slv13_arvalid(slv13_arvalid)
    ,.slv13_awaddr(slv13_awaddr[31:0])
    ,.slv13_awburst(slv13_awburst[1:0])
    ,.slv13_awextras(slv13_awextras[(EXTRAS - 1):0])
    ,.slv13_awid(slv13_awid[(IDWID - 1):0])
    ,.slv13_awlen(slv13_awlen[7:0])
    ,.slv13_awready(slv13_awready)
    ,.slv13_awvalid(slv13_awvalid)
    ,.slv13_bid(slv13_bid[(IDWID - 1):0])
    ,.slv13_bready(slv13_bready)
    ,.slv13_bresp(slv13_bresp[1:0])
    ,.slv13_bvalid(slv13_bvalid)
    ,.slv13_rdata(slv13_rdata[(DWID - 1):0])
    ,.slv13_rid(slv13_rid[(IDWID - 1):0])
    ,.slv13_rlast(slv13_rlast)
    ,.slv13_rready(slv13_rready)
    ,.slv13_rresp(slv13_rresp[1:0])
    ,.slv13_rvalid(slv13_rvalid)
    ,.slv13_wdata(slv13_wdata[(DWID - 1):0])
    ,.slv13_wlast(slv13_wlast)
    ,.slv13_wready(slv13_wready)
    ,.slv13_wstrb(slv13_wstrb[(WSTRB - 1):0])
    ,.slv13_wvalid(slv13_wvalid)


    ,.slv14_araddr(slv14_araddr[31:0])
    ,.slv14_arburst(slv14_arburst[1:0])
    ,.slv14_arextras(slv14_arextras[(EXTRAS - 1):0])
    ,.slv14_arid(slv14_arid[(IDWID - 1):0])
    ,.slv14_arlen(slv14_arlen[7:0])
    ,.slv14_arready(slv14_arready)
    ,.slv14_arvalid(slv14_arvalid)
    ,.slv14_awaddr(slv14_awaddr[31:0])
    ,.slv14_awburst(slv14_awburst[1:0])
    ,.slv14_awextras(slv14_awextras[(EXTRAS - 1):0])
    ,.slv14_awid(slv14_awid[(IDWID - 1):0])
    ,.slv14_awlen(slv14_awlen[7:0])
    ,.slv14_awready(slv14_awready)
    ,.slv14_awvalid(slv14_awvalid)
    ,.slv14_bid(slv14_bid[(IDWID - 1):0])
    ,.slv14_bready(slv14_bready)
    ,.slv14_bresp(slv14_bresp[1:0])
    ,.slv14_bvalid(slv14_bvalid)
    ,.slv14_rdata(slv14_rdata[(DWID - 1):0])
    ,.slv14_rid(slv14_rid[(IDWID - 1):0])
    ,.slv14_rlast(slv14_rlast)
    ,.slv14_rready(slv14_rready)
    ,.slv14_rresp(slv14_rresp[1:0])
    ,.slv14_rvalid(slv14_rvalid)
    ,.slv14_wdata(slv14_wdata[(DWID - 1):0])
    ,.slv14_wlast(slv14_wlast)
    ,.slv14_wready(slv14_wready)
    ,.slv14_wstrb(slv14_wstrb[(WSTRB - 1):0])
    ,.slv14_wvalid(slv14_wvalid)


    ,.slv15_araddr(slv15_araddr[31:0])
    ,.slv15_arburst(slv15_arburst[1:0])
    ,.slv15_arextras(slv15_arextras[(EXTRAS - 1):0])
    ,.slv15_arid(slv15_arid[(IDWID - 1):0])
    ,.slv15_arlen(slv15_arlen[7:0])
    ,.slv15_arready(slv15_arready)
    ,.slv15_arvalid(slv15_arvalid)
    ,.slv15_awaddr(slv15_awaddr[31:0])
    ,.slv15_awburst(slv15_awburst[1:0])
    ,.slv15_awextras(slv15_awextras[(EXTRAS - 1):0])
    ,.slv15_awid(slv15_awid[(IDWID - 1):0])
    ,.slv15_awlen(slv15_awlen[7:0])
    ,.slv15_awready(slv15_awready)
    ,.slv15_awvalid(slv15_awvalid)
    ,.slv15_bid(slv15_bid[(IDWID - 1):0])
    ,.slv15_bready(slv15_bready)
    ,.slv15_bresp(slv15_bresp[1:0])
    ,.slv15_bvalid(slv15_bvalid)
    ,.slv15_rdata(slv15_rdata[(DWID - 1):0])
    ,.slv15_rid(slv15_rid[(IDWID - 1):0])
    ,.slv15_rlast(slv15_rlast)
    ,.slv15_rready(slv15_rready)
    ,.slv15_rresp(slv15_rresp[1:0])
    ,.slv15_rvalid(slv15_rvalid)
    ,.slv15_wdata(slv15_wdata[(DWID - 1):0])
    ,.slv15_wlast(slv15_wlast)
    ,.slv15_wready(slv15_wready)
    ,.slv15_wstrb(slv15_wstrb[(WSTRB - 1):0])
    ,.slv15_wvalid(slv15_wvalid)


    ,.slv2_araddr(slv2_araddr[31:0])
    ,.slv2_arburst(slv2_arburst[1:0])
    ,.slv2_arextras(slv2_arextras[(EXTRAS - 1):0])
    ,.slv2_arid(slv2_arid[(IDWID - 1):0])
    ,.slv2_arlen(slv2_arlen[7:0])
    ,.slv2_arready(slv2_arready)
    ,.slv2_arvalid(slv2_arvalid)
    ,.slv2_awaddr(slv2_awaddr[31:0])
    ,.slv2_awburst(slv2_awburst[1:0])
    ,.slv2_awextras(slv2_awextras[(EXTRAS - 1):0])
    ,.slv2_awid(slv2_awid[(IDWID - 1):0])
    ,.slv2_awlen(slv2_awlen[7:0])
    ,.slv2_awready(slv2_awready)
    ,.slv2_awvalid(slv2_awvalid)
    ,.slv2_bid(slv2_bid[(IDWID - 1):0])
    ,.slv2_bready(slv2_bready)
    ,.slv2_bresp(slv2_bresp[1:0])
    ,.slv2_bvalid(slv2_bvalid)
    ,.slv2_rdata(slv2_rdata[(DWID - 1):0])
    ,.slv2_rid(slv2_rid[(IDWID - 1):0])
    ,.slv2_rlast(slv2_rlast)
    ,.slv2_rready(slv2_rready)
    ,.slv2_rresp(slv2_rresp[1:0])
    ,.slv2_rvalid(slv2_rvalid)
    ,.slv2_wdata(slv2_wdata[(DWID - 1):0])
    ,.slv2_wlast(slv2_wlast)
    ,.slv2_wready(slv2_wready)
    ,.slv2_wstrb(slv2_wstrb[(WSTRB - 1):0])
    ,.slv2_wvalid(slv2_wvalid)


    ,.slv3_araddr(slv3_araddr[31:0])
    ,.slv3_arburst(slv3_arburst[1:0])
    ,.slv3_arextras(slv3_arextras[(EXTRAS - 1):0])
    ,.slv3_arid(slv3_arid[(IDWID - 1):0])
    ,.slv3_arlen(slv3_arlen[7:0])
    ,.slv3_arready(slv3_arready)
    ,.slv3_arvalid(slv3_arvalid)
    ,.slv3_awaddr(slv3_awaddr[31:0])
    ,.slv3_awburst(slv3_awburst[1:0])
    ,.slv3_awextras(slv3_awextras[(EXTRAS - 1):0])
    ,.slv3_awid(slv3_awid[(IDWID - 1):0])
    ,.slv3_awlen(slv3_awlen[7:0])
    ,.slv3_awready(slv3_awready)
    ,.slv3_awvalid(slv3_awvalid)
    ,.slv3_bid(slv3_bid[(IDWID - 1):0])
    ,.slv3_bready(slv3_bready)
    ,.slv3_bresp(slv3_bresp[1:0])
    ,.slv3_bvalid(slv3_bvalid)
    ,.slv3_rdata(slv3_rdata[(DWID - 1):0])
    ,.slv3_rid(slv3_rid[(IDWID - 1):0])
    ,.slv3_rlast(slv3_rlast)
    ,.slv3_rready(slv3_rready)
    ,.slv3_rresp(slv3_rresp[1:0])
    ,.slv3_rvalid(slv3_rvalid)
    ,.slv3_wdata(slv3_wdata[(DWID - 1):0])
    ,.slv3_wlast(slv3_wlast)
    ,.slv3_wready(slv3_wready)
    ,.slv3_wstrb(slv3_wstrb[(WSTRB - 1):0])
    ,.slv3_wvalid(slv3_wvalid)


    ,.slv4_araddr(slv4_araddr[31:0])
    ,.slv4_arburst(slv4_arburst[1:0])
    ,.slv4_arextras(slv4_arextras[(EXTRAS - 1):0])
    ,.slv4_arid(slv4_arid[(IDWID - 1):0])
    ,.slv4_arlen(slv4_arlen[7:0])
    ,.slv4_arready(slv4_arready)
    ,.slv4_arvalid(slv4_arvalid)
    ,.slv4_awaddr(slv4_awaddr[31:0])
    ,.slv4_awburst(slv4_awburst[1:0])
    ,.slv4_awextras(slv4_awextras[(EXTRAS - 1):0])
    ,.slv4_awid(slv4_awid[(IDWID - 1):0])
    ,.slv4_awlen(slv4_awlen[7:0])
    ,.slv4_awready(slv4_awready)
    ,.slv4_awvalid(slv4_awvalid)
    ,.slv4_bid(slv4_bid[(IDWID - 1):0])
    ,.slv4_bready(slv4_bready)
    ,.slv4_bresp(slv4_bresp[1:0])
    ,.slv4_bvalid(slv4_bvalid)
    ,.slv4_rdata(slv4_rdata[(DWID - 1):0])
    ,.slv4_rid(slv4_rid[(IDWID - 1):0])
    ,.slv4_rlast(slv4_rlast)
    ,.slv4_rready(slv4_rready)
    ,.slv4_rresp(slv4_rresp[1:0])
    ,.slv4_rvalid(slv4_rvalid)
    ,.slv4_wdata(slv4_wdata[(DWID - 1):0])
    ,.slv4_wlast(slv4_wlast)
    ,.slv4_wready(slv4_wready)
    ,.slv4_wstrb(slv4_wstrb[(WSTRB - 1):0])
    ,.slv4_wvalid(slv4_wvalid)


    ,.slv5_araddr(slv5_araddr[31:0])
    ,.slv5_arburst(slv5_arburst[1:0])
    ,.slv5_arextras(slv5_arextras[(EXTRAS - 1):0])
    ,.slv5_arid(slv5_arid[(IDWID - 1):0])
    ,.slv5_arlen(slv5_arlen[7:0])
    ,.slv5_arready(slv5_arready)
    ,.slv5_arvalid(slv5_arvalid)
    ,.slv5_awaddr(slv5_awaddr[31:0])
    ,.slv5_awburst(slv5_awburst[1:0])
    ,.slv5_awextras(slv5_awextras[(EXTRAS - 1):0])
    ,.slv5_awid(slv5_awid[(IDWID - 1):0])
    ,.slv5_awlen(slv5_awlen[7:0])
    ,.slv5_awready(slv5_awready)
    ,.slv5_awvalid(slv5_awvalid)
    ,.slv5_bid(slv5_bid[(IDWID - 1):0])
    ,.slv5_bready(slv5_bready)
    ,.slv5_bresp(slv5_bresp[1:0])
    ,.slv5_bvalid(slv5_bvalid)
    ,.slv5_rdata(slv5_rdata[(DWID - 1):0])
    ,.slv5_rid(slv5_rid[(IDWID - 1):0])
    ,.slv5_rlast(slv5_rlast)
    ,.slv5_rready(slv5_rready)
    ,.slv5_rresp(slv5_rresp[1:0])
    ,.slv5_rvalid(slv5_rvalid)
    ,.slv5_wdata(slv5_wdata[(DWID - 1):0])
    ,.slv5_wlast(slv5_wlast)
    ,.slv5_wready(slv5_wready)
    ,.slv5_wstrb(slv5_wstrb[(WSTRB - 1):0])
    ,.slv5_wvalid(slv5_wvalid)


    ,.slv6_araddr(slv6_araddr[31:0])
    ,.slv6_arburst(slv6_arburst[1:0])
    ,.slv6_arextras(slv6_arextras[(EXTRAS - 1):0])
    ,.slv6_arid(slv6_arid[(IDWID - 1):0])
    ,.slv6_arlen(slv6_arlen[7:0])
    ,.slv6_arready(slv6_arready)
    ,.slv6_arvalid(slv6_arvalid)
    ,.slv6_awaddr(slv6_awaddr[31:0])
    ,.slv6_awburst(slv6_awburst[1:0])
    ,.slv6_awextras(slv6_awextras[(EXTRAS - 1):0])
    ,.slv6_awid(slv6_awid[(IDWID - 1):0])
    ,.slv6_awlen(slv6_awlen[7:0])
    ,.slv6_awready(slv6_awready)
    ,.slv6_awvalid(slv6_awvalid)
    ,.slv6_bid(slv6_bid[(IDWID - 1):0])
    ,.slv6_bready(slv6_bready)
    ,.slv6_bresp(slv6_bresp[1:0])
    ,.slv6_bvalid(slv6_bvalid)
    ,.slv6_rdata(slv6_rdata[(DWID - 1):0])
    ,.slv6_rid(slv6_rid[(IDWID - 1):0])
    ,.slv6_rlast(slv6_rlast)
    ,.slv6_rready(slv6_rready)
    ,.slv6_rresp(slv6_rresp[1:0])
    ,.slv6_rvalid(slv6_rvalid)
    ,.slv6_wdata(slv6_wdata[(DWID - 1):0])
    ,.slv6_wlast(slv6_wlast)
    ,.slv6_wready(slv6_wready)
    ,.slv6_wstrb(slv6_wstrb[(WSTRB - 1):0])
    ,.slv6_wvalid(slv6_wvalid)


    ,.slv7_araddr(slv7_araddr[31:0])
    ,.slv7_arburst(slv7_arburst[1:0])
    ,.slv7_arextras(slv7_arextras[(EXTRAS - 1):0])
    ,.slv7_arid(slv7_arid[(IDWID - 1):0])
    ,.slv7_arlen(slv7_arlen[7:0])
    ,.slv7_arready(slv7_arready)
    ,.slv7_arvalid(slv7_arvalid)
    ,.slv7_awaddr(slv7_awaddr[31:0])
    ,.slv7_awburst(slv7_awburst[1:0])
    ,.slv7_awextras(slv7_awextras[(EXTRAS - 1):0])
    ,.slv7_awid(slv7_awid[(IDWID - 1):0])
    ,.slv7_awlen(slv7_awlen[7:0])
    ,.slv7_awready(slv7_awready)
    ,.slv7_awvalid(slv7_awvalid)
    ,.slv7_bid(slv7_bid[(IDWID - 1):0])
    ,.slv7_bready(slv7_bready)
    ,.slv7_bresp(slv7_bresp[1:0])
    ,.slv7_bvalid(slv7_bvalid)
    ,.slv7_rdata(slv7_rdata[(DWID - 1):0])
    ,.slv7_rid(slv7_rid[(IDWID - 1):0])
    ,.slv7_rlast(slv7_rlast)
    ,.slv7_rready(slv7_rready)
    ,.slv7_rresp(slv7_rresp[1:0])
    ,.slv7_rvalid(slv7_rvalid)
    ,.slv7_wdata(slv7_wdata[(DWID - 1):0])
    ,.slv7_wlast(slv7_wlast)
    ,.slv7_wready(slv7_wready)
    ,.slv7_wstrb(slv7_wstrb[(WSTRB - 1):0])
    ,.slv7_wvalid(slv7_wvalid)


    ,.slv8_araddr(slv8_araddr[31:0])
    ,.slv8_arburst(slv8_arburst[1:0])
    ,.slv8_arextras(slv8_arextras[(EXTRAS - 1):0])
    ,.slv8_arid(slv8_arid[(IDWID - 1):0])
    ,.slv8_arlen(slv8_arlen[7:0])
    ,.slv8_arready(slv8_arready)
    ,.slv8_arvalid(slv8_arvalid)
    ,.slv8_awaddr(slv8_awaddr[31:0])
    ,.slv8_awburst(slv8_awburst[1:0])
    ,.slv8_awextras(slv8_awextras[(EXTRAS - 1):0])
    ,.slv8_awid(slv8_awid[(IDWID - 1):0])
    ,.slv8_awlen(slv8_awlen[7:0])
    ,.slv8_awready(slv8_awready)
    ,.slv8_awvalid(slv8_awvalid)
    ,.slv8_bid(slv8_bid[(IDWID - 1):0])
    ,.slv8_bready(slv8_bready)
    ,.slv8_bresp(slv8_bresp[1:0])
    ,.slv8_bvalid(slv8_bvalid)
    ,.slv8_rdata(slv8_rdata[(DWID - 1):0])
    ,.slv8_rid(slv8_rid[(IDWID - 1):0])
    ,.slv8_rlast(slv8_rlast)
    ,.slv8_rready(slv8_rready)
    ,.slv8_rresp(slv8_rresp[1:0])
    ,.slv8_rvalid(slv8_rvalid)
    ,.slv8_wdata(slv8_wdata[(DWID - 1):0])
    ,.slv8_wlast(slv8_wlast)
    ,.slv8_wready(slv8_wready)
    ,.slv8_wstrb(slv8_wstrb[(WSTRB - 1):0])
    ,.slv8_wvalid(slv8_wvalid)


    ,.slv9_araddr(slv9_araddr[31:0])
    ,.slv9_arburst(slv9_arburst[1:0])
    ,.slv9_arextras(slv9_arextras[(EXTRAS - 1):0])
    ,.slv9_arid(slv9_arid[(IDWID - 1):0])
    ,.slv9_arlen(slv9_arlen[7:0])
    ,.slv9_arready(slv9_arready)
    ,.slv9_arvalid(slv9_arvalid)
    ,.slv9_awaddr(slv9_awaddr[31:0])
    ,.slv9_awburst(slv9_awburst[1:0])
    ,.slv9_awextras(slv9_awextras[(EXTRAS - 1):0])
    ,.slv9_awid(slv9_awid[(IDWID - 1):0])
    ,.slv9_awlen(slv9_awlen[7:0])
    ,.slv9_awready(slv9_awready)
    ,.slv9_awvalid(slv9_awvalid)
    ,.slv9_bid(slv9_bid[(IDWID - 1):0])
    ,.slv9_bready(slv9_bready)
    ,.slv9_bresp(slv9_bresp[1:0])
    ,.slv9_bvalid(slv9_bvalid)
    ,.slv9_rdata(slv9_rdata[(DWID - 1):0])
    ,.slv9_rid(slv9_rid[(IDWID - 1):0])
    ,.slv9_rlast(slv9_rlast)
    ,.slv9_rready(slv9_rready)
    ,.slv9_rresp(slv9_rresp[1:0])
    ,.slv9_rvalid(slv9_rvalid)
    ,.slv9_wdata(slv9_wdata[(DWID - 1):0])
    ,.slv9_wlast(slv9_wlast)
    ,.slv9_wready(slv9_wready)
    ,.slv9_wstrb(slv9_wstrb[(WSTRB - 1):0])
    ,.slv9_wvalid(slv9_wvalid)


    ,.mst0_araddr(mst0_araddr[31:0])
    ,.mst0_arburst(mst0_arburst[1:0])
    ,.mst0_arextras(mst0_arextras[(EXTRAS - 1):0])
    ,.mst0_arid(mst0_arid[(IDWID - 1):0])
    ,.mst0_arlen(mst0_arlen[7:0])
    ,.mst0_arready(mst0_arready)
    ,.mst0_arvalid(mst0_arvalid)
    ,.mst0_awaddr(mst0_awaddr[31:0])
    ,.mst0_awburst(mst0_awburst[1:0])
    ,.mst0_awextras(mst0_awextras[(EXTRAS - 1):0])
    ,.mst0_awid(mst0_awid[(IDWID - 1):0])
    ,.mst0_awlen(mst0_awlen[7:0])
    ,.mst0_awready(mst0_awready)
    ,.mst0_awvalid(mst0_awvalid)
    ,.mst0_bid(mst0_bid[(IDWID - 1):0])
    ,.mst0_bready(mst0_bready)
    ,.mst0_bresp(mst0_bresp[1:0])
    ,.mst0_bvalid(mst0_bvalid)
    ,.mst0_rdata(mst0_rdata[(DWID - 1):0])
    ,.mst0_rid(mst0_rid[(IDWID - 1):0])
    ,.mst0_rlast(mst0_rlast)
    ,.mst0_rready(mst0_rready)
    ,.mst0_rresp(mst0_rresp[1:0])
    ,.mst0_rvalid(mst0_rvalid)
    ,.mst0_wdata(mst0_wdata[(DWID - 1):0])
    ,.mst0_wlast(mst0_wlast)
    ,.mst0_wready(mst0_wready)
    ,.mst0_wstrb(mst0_wstrb[(WSTRB - 1):0])
    ,.mst0_wvalid(mst0_wvalid)

    ,.mst1_araddr(mst1_araddr[31:0])
    ,.mst1_arburst(mst1_arburst[1:0])
    ,.mst1_arextras(mst1_arextras[(EXTRAS - 1):0])
    ,.mst1_arid(mst1_arid[(IDWID - 1):0])
    ,.mst1_arlen(mst1_arlen[7:0])
    ,.mst1_arready(mst1_arready)
    ,.mst1_arvalid(mst1_arvalid)
    ,.mst1_awaddr(mst1_awaddr[31:0])
    ,.mst1_awburst(mst1_awburst[1:0])
    ,.mst1_awextras(mst1_awextras[(EXTRAS - 1):0])
    ,.mst1_awid(mst1_awid[(IDWID - 1):0])
    ,.mst1_awlen(mst1_awlen[7:0])
    ,.mst1_awready(mst1_awready)
    ,.mst1_awvalid(mst1_awvalid)
    ,.mst1_bid(mst1_bid[(IDWID - 1):0])
    ,.mst1_bready(mst1_bready)
    ,.mst1_bresp(mst1_bresp[1:0])
    ,.mst1_bvalid(mst1_bvalid)
    ,.mst1_rdata(mst1_rdata[(DWID - 1):0])
    ,.mst1_rid(mst1_rid[(IDWID - 1):0])
    ,.mst1_rlast(mst1_rlast)
    ,.mst1_rready(mst1_rready)
    ,.mst1_rresp(mst1_rresp[1:0])
    ,.mst1_rvalid(mst1_rvalid)
    ,.mst1_wdata(mst1_wdata[(DWID - 1):0])
    ,.mst1_wlast(mst1_wlast)
    ,.mst1_wready(mst1_wready)
    ,.mst1_wstrb(mst1_wstrb[(WSTRB - 1):0])
    ,.mst1_wvalid(mst1_wvalid)

    ,.mst10_araddr(mst10_araddr[31:0])
    ,.mst10_arburst(mst10_arburst[1:0])
    ,.mst10_arextras(mst10_arextras[(EXTRAS - 1):0])
    ,.mst10_arid(mst10_arid[(IDWID - 1):0])
    ,.mst10_arlen(mst10_arlen[7:0])
    ,.mst10_arready(mst10_arready)
    ,.mst10_arvalid(mst10_arvalid)
    ,.mst10_awaddr(mst10_awaddr[31:0])
    ,.mst10_awburst(mst10_awburst[1:0])
    ,.mst10_awextras(mst10_awextras[(EXTRAS - 1):0])
    ,.mst10_awid(mst10_awid[(IDWID - 1):0])
    ,.mst10_awlen(mst10_awlen[7:0])
    ,.mst10_awready(mst10_awready)
    ,.mst10_awvalid(mst10_awvalid)
    ,.mst10_bid(mst10_bid[(IDWID - 1):0])
    ,.mst10_bready(mst10_bready)
    ,.mst10_bresp(mst10_bresp[1:0])
    ,.mst10_bvalid(mst10_bvalid)
    ,.mst10_rdata(mst10_rdata[(DWID - 1):0])
    ,.mst10_rid(mst10_rid[(IDWID - 1):0])
    ,.mst10_rlast(mst10_rlast)
    ,.mst10_rready(mst10_rready)
    ,.mst10_rresp(mst10_rresp[1:0])
    ,.mst10_rvalid(mst10_rvalid)
    ,.mst10_wdata(mst10_wdata[(DWID - 1):0])
    ,.mst10_wlast(mst10_wlast)
    ,.mst10_wready(mst10_wready)
    ,.mst10_wstrb(mst10_wstrb[(WSTRB - 1):0])
    ,.mst10_wvalid(mst10_wvalid)

    ,.mst11_araddr(mst11_araddr[31:0])
    ,.mst11_arburst(mst11_arburst[1:0])
    ,.mst11_arextras(mst11_arextras[(EXTRAS - 1):0])
    ,.mst11_arid(mst11_arid[(IDWID - 1):0])
    ,.mst11_arlen(mst11_arlen[7:0])
    ,.mst11_arready(mst11_arready)
    ,.mst11_arvalid(mst11_arvalid)
    ,.mst11_awaddr(mst11_awaddr[31:0])
    ,.mst11_awburst(mst11_awburst[1:0])
    ,.mst11_awextras(mst11_awextras[(EXTRAS - 1):0])
    ,.mst11_awid(mst11_awid[(IDWID - 1):0])
    ,.mst11_awlen(mst11_awlen[7:0])
    ,.mst11_awready(mst11_awready)
    ,.mst11_awvalid(mst11_awvalid)
    ,.mst11_bid(mst11_bid[(IDWID - 1):0])
    ,.mst11_bready(mst11_bready)
    ,.mst11_bresp(mst11_bresp[1:0])
    ,.mst11_bvalid(mst11_bvalid)
    ,.mst11_rdata(mst11_rdata[(DWID - 1):0])
    ,.mst11_rid(mst11_rid[(IDWID - 1):0])
    ,.mst11_rlast(mst11_rlast)
    ,.mst11_rready(mst11_rready)
    ,.mst11_rresp(mst11_rresp[1:0])
    ,.mst11_rvalid(mst11_rvalid)
    ,.mst11_wdata(mst11_wdata[(DWID - 1):0])
    ,.mst11_wlast(mst11_wlast)
    ,.mst11_wready(mst11_wready)
    ,.mst11_wstrb(mst11_wstrb[(WSTRB - 1):0])
    ,.mst11_wvalid(mst11_wvalid)

    ,.mst12_araddr(mst12_araddr[31:0])
    ,.mst12_arburst(mst12_arburst[1:0])
    ,.mst12_arextras(mst12_arextras[(EXTRAS - 1):0])
    ,.mst12_arid(mst12_arid[(IDWID - 1):0])
    ,.mst12_arlen(mst12_arlen[7:0])
    ,.mst12_arready(mst12_arready)
    ,.mst12_arvalid(mst12_arvalid)
    ,.mst12_awaddr(mst12_awaddr[31:0])
    ,.mst12_awburst(mst12_awburst[1:0])
    ,.mst12_awextras(mst12_awextras[(EXTRAS - 1):0])
    ,.mst12_awid(mst12_awid[(IDWID - 1):0])
    ,.mst12_awlen(mst12_awlen[7:0])
    ,.mst12_awready(mst12_awready)
    ,.mst12_awvalid(mst12_awvalid)
    ,.mst12_bid(mst12_bid[(IDWID - 1):0])
    ,.mst12_bready(mst12_bready)
    ,.mst12_bresp(mst12_bresp[1:0])
    ,.mst12_bvalid(mst12_bvalid)
    ,.mst12_rdata(mst12_rdata[(DWID - 1):0])
    ,.mst12_rid(mst12_rid[(IDWID - 1):0])
    ,.mst12_rlast(mst12_rlast)
    ,.mst12_rready(mst12_rready)
    ,.mst12_rresp(mst12_rresp[1:0])
    ,.mst12_rvalid(mst12_rvalid)
    ,.mst12_wdata(mst12_wdata[(DWID - 1):0])
    ,.mst12_wlast(mst12_wlast)
    ,.mst12_wready(mst12_wready)
    ,.mst12_wstrb(mst12_wstrb[(WSTRB - 1):0])
    ,.mst12_wvalid(mst12_wvalid)

    ,.mst13_araddr(mst13_araddr[31:0])
    ,.mst13_arburst(mst13_arburst[1:0])
    ,.mst13_arextras(mst13_arextras[(EXTRAS - 1):0])
    ,.mst13_arid(mst13_arid[(IDWID - 1):0])
    ,.mst13_arlen(mst13_arlen[7:0])
    ,.mst13_arready(mst13_arready)
    ,.mst13_arvalid(mst13_arvalid)
    ,.mst13_awaddr(mst13_awaddr[31:0])
    ,.mst13_awburst(mst13_awburst[1:0])
    ,.mst13_awextras(mst13_awextras[(EXTRAS - 1):0])
    ,.mst13_awid(mst13_awid[(IDWID - 1):0])
    ,.mst13_awlen(mst13_awlen[7:0])
    ,.mst13_awready(mst13_awready)
    ,.mst13_awvalid(mst13_awvalid)
    ,.mst13_bid(mst13_bid[(IDWID - 1):0])
    ,.mst13_bready(mst13_bready)
    ,.mst13_bresp(mst13_bresp[1:0])
    ,.mst13_bvalid(mst13_bvalid)
    ,.mst13_rdata(mst13_rdata[(DWID - 1):0])
    ,.mst13_rid(mst13_rid[(IDWID - 1):0])
    ,.mst13_rlast(mst13_rlast)
    ,.mst13_rready(mst13_rready)
    ,.mst13_rresp(mst13_rresp[1:0])
    ,.mst13_rvalid(mst13_rvalid)
    ,.mst13_wdata(mst13_wdata[(DWID - 1):0])
    ,.mst13_wlast(mst13_wlast)
    ,.mst13_wready(mst13_wready)
    ,.mst13_wstrb(mst13_wstrb[(WSTRB - 1):0])
    ,.mst13_wvalid(mst13_wvalid)

    ,.mst14_araddr(mst14_araddr[31:0])
    ,.mst14_arburst(mst14_arburst[1:0])
    ,.mst14_arextras(mst14_arextras[(EXTRAS - 1):0])
    ,.mst14_arid(mst14_arid[(IDWID - 1):0])
    ,.mst14_arlen(mst14_arlen[7:0])
    ,.mst14_arready(mst14_arready)
    ,.mst14_arvalid(mst14_arvalid)
    ,.mst14_awaddr(mst14_awaddr[31:0])
    ,.mst14_awburst(mst14_awburst[1:0])
    ,.mst14_awextras(mst14_awextras[(EXTRAS - 1):0])
    ,.mst14_awid(mst14_awid[(IDWID - 1):0])
    ,.mst14_awlen(mst14_awlen[7:0])
    ,.mst14_awready(mst14_awready)
    ,.mst14_awvalid(mst14_awvalid)
    ,.mst14_bid(mst14_bid[(IDWID - 1):0])
    ,.mst14_bready(mst14_bready)
    ,.mst14_bresp(mst14_bresp[1:0])
    ,.mst14_bvalid(mst14_bvalid)
    ,.mst14_rdata(mst14_rdata[(DWID - 1):0])
    ,.mst14_rid(mst14_rid[(IDWID - 1):0])
    ,.mst14_rlast(mst14_rlast)
    ,.mst14_rready(mst14_rready)
    ,.mst14_rresp(mst14_rresp[1:0])
    ,.mst14_rvalid(mst14_rvalid)
    ,.mst14_wdata(mst14_wdata[(DWID - 1):0])
    ,.mst14_wlast(mst14_wlast)
    ,.mst14_wready(mst14_wready)
    ,.mst14_wstrb(mst14_wstrb[(WSTRB - 1):0])
    ,.mst14_wvalid(mst14_wvalid)

    ,.mst15_araddr(mst15_araddr[31:0])
    ,.mst15_arburst(mst15_arburst[1:0])
    ,.mst15_arextras(mst15_arextras[(EXTRAS - 1):0])
    ,.mst15_arid(mst15_arid[(IDWID - 1):0])
    ,.mst15_arlen(mst15_arlen[7:0])
    ,.mst15_arready(mst15_arready)
    ,.mst15_arvalid(mst15_arvalid)
    ,.mst15_awaddr(mst15_awaddr[31:0])
    ,.mst15_awburst(mst15_awburst[1:0])
    ,.mst15_awextras(mst15_awextras[(EXTRAS - 1):0])
    ,.mst15_awid(mst15_awid[(IDWID - 1):0])
    ,.mst15_awlen(mst15_awlen[7:0])
    ,.mst15_awready(mst15_awready)
    ,.mst15_awvalid(mst15_awvalid)
    ,.mst15_bid(mst15_bid[(IDWID - 1):0])
    ,.mst15_bready(mst15_bready)
    ,.mst15_bresp(mst15_bresp[1:0])
    ,.mst15_bvalid(mst15_bvalid)
    ,.mst15_rdata(mst15_rdata[(DWID - 1):0])
    ,.mst15_rid(mst15_rid[(IDWID - 1):0])
    ,.mst15_rlast(mst15_rlast)
    ,.mst15_rready(mst15_rready)
    ,.mst15_rresp(mst15_rresp[1:0])
    ,.mst15_rvalid(mst15_rvalid)
    ,.mst15_wdata(mst15_wdata[(DWID - 1):0])
    ,.mst15_wlast(mst15_wlast)
    ,.mst15_wready(mst15_wready)
    ,.mst15_wstrb(mst15_wstrb[(WSTRB - 1):0])
    ,.mst15_wvalid(mst15_wvalid)

    ,.mst2_araddr(mst2_araddr[31:0])
    ,.mst2_arburst(mst2_arburst[1:0])
    ,.mst2_arextras(mst2_arextras[(EXTRAS - 1):0])
    ,.mst2_arid(mst2_arid[(IDWID - 1):0])
    ,.mst2_arlen(mst2_arlen[7:0])
    ,.mst2_arready(mst2_arready)
    ,.mst2_arvalid(mst2_arvalid)
    ,.mst2_awaddr(mst2_awaddr[31:0])
    ,.mst2_awburst(mst2_awburst[1:0])
    ,.mst2_awextras(mst2_awextras[(EXTRAS - 1):0])
    ,.mst2_awid(mst2_awid[(IDWID - 1):0])
    ,.mst2_awlen(mst2_awlen[7:0])
    ,.mst2_awready(mst2_awready)
    ,.mst2_awvalid(mst2_awvalid)
    ,.mst2_bid(mst2_bid[(IDWID - 1):0])
    ,.mst2_bready(mst2_bready)
    ,.mst2_bresp(mst2_bresp[1:0])
    ,.mst2_bvalid(mst2_bvalid)
    ,.mst2_rdata(mst2_rdata[(DWID - 1):0])
    ,.mst2_rid(mst2_rid[(IDWID - 1):0])
    ,.mst2_rlast(mst2_rlast)
    ,.mst2_rready(mst2_rready)
    ,.mst2_rresp(mst2_rresp[1:0])
    ,.mst2_rvalid(mst2_rvalid)
    ,.mst2_wdata(mst2_wdata[(DWID - 1):0])
    ,.mst2_wlast(mst2_wlast)
    ,.mst2_wready(mst2_wready)
    ,.mst2_wstrb(mst2_wstrb[(WSTRB - 1):0])
    ,.mst2_wvalid(mst2_wvalid)

    ,.mst3_araddr(mst3_araddr[31:0])
    ,.mst3_arburst(mst3_arburst[1:0])
    ,.mst3_arextras(mst3_arextras[(EXTRAS - 1):0])
    ,.mst3_arid(mst3_arid[(IDWID - 1):0])
    ,.mst3_arlen(mst3_arlen[7:0])
    ,.mst3_arready(mst3_arready)
    ,.mst3_arvalid(mst3_arvalid)
    ,.mst3_awaddr(mst3_awaddr[31:0])
    ,.mst3_awburst(mst3_awburst[1:0])
    ,.mst3_awextras(mst3_awextras[(EXTRAS - 1):0])
    ,.mst3_awid(mst3_awid[(IDWID - 1):0])
    ,.mst3_awlen(mst3_awlen[7:0])
    ,.mst3_awready(mst3_awready)
    ,.mst3_awvalid(mst3_awvalid)
    ,.mst3_bid(mst3_bid[(IDWID - 1):0])
    ,.mst3_bready(mst3_bready)
    ,.mst3_bresp(mst3_bresp[1:0])
    ,.mst3_bvalid(mst3_bvalid)
    ,.mst3_rdata(mst3_rdata[(DWID - 1):0])
    ,.mst3_rid(mst3_rid[(IDWID - 1):0])
    ,.mst3_rlast(mst3_rlast)
    ,.mst3_rready(mst3_rready)
    ,.mst3_rresp(mst3_rresp[1:0])
    ,.mst3_rvalid(mst3_rvalid)
    ,.mst3_wdata(mst3_wdata[(DWID - 1):0])
    ,.mst3_wlast(mst3_wlast)
    ,.mst3_wready(mst3_wready)
    ,.mst3_wstrb(mst3_wstrb[(WSTRB - 1):0])
    ,.mst3_wvalid(mst3_wvalid)

    ,.mst4_araddr(mst4_araddr[31:0])
    ,.mst4_arburst(mst4_arburst[1:0])
    ,.mst4_arextras(mst4_arextras[(EXTRAS - 1):0])
    ,.mst4_arid(mst4_arid[(IDWID - 1):0])
    ,.mst4_arlen(mst4_arlen[7:0])
    ,.mst4_arready(mst4_arready)
    ,.mst4_arvalid(mst4_arvalid)
    ,.mst4_awaddr(mst4_awaddr[31:0])
    ,.mst4_awburst(mst4_awburst[1:0])
    ,.mst4_awextras(mst4_awextras[(EXTRAS - 1):0])
    ,.mst4_awid(mst4_awid[(IDWID - 1):0])
    ,.mst4_awlen(mst4_awlen[7:0])
    ,.mst4_awready(mst4_awready)
    ,.mst4_awvalid(mst4_awvalid)
    ,.mst4_bid(mst4_bid[(IDWID - 1):0])
    ,.mst4_bready(mst4_bready)
    ,.mst4_bresp(mst4_bresp[1:0])
    ,.mst4_bvalid(mst4_bvalid)
    ,.mst4_rdata(mst4_rdata[(DWID - 1):0])
    ,.mst4_rid(mst4_rid[(IDWID - 1):0])
    ,.mst4_rlast(mst4_rlast)
    ,.mst4_rready(mst4_rready)
    ,.mst4_rresp(mst4_rresp[1:0])
    ,.mst4_rvalid(mst4_rvalid)
    ,.mst4_wdata(mst4_wdata[(DWID - 1):0])
    ,.mst4_wlast(mst4_wlast)
    ,.mst4_wready(mst4_wready)
    ,.mst4_wstrb(mst4_wstrb[(WSTRB - 1):0])
    ,.mst4_wvalid(mst4_wvalid)

    ,.mst5_araddr(mst5_araddr[31:0])
    ,.mst5_arburst(mst5_arburst[1:0])
    ,.mst5_arextras(mst5_arextras[(EXTRAS - 1):0])
    ,.mst5_arid(mst5_arid[(IDWID - 1):0])
    ,.mst5_arlen(mst5_arlen[7:0])
    ,.mst5_arready(mst5_arready)
    ,.mst5_arvalid(mst5_arvalid)
    ,.mst5_awaddr(mst5_awaddr[31:0])
    ,.mst5_awburst(mst5_awburst[1:0])
    ,.mst5_awextras(mst5_awextras[(EXTRAS - 1):0])
    ,.mst5_awid(mst5_awid[(IDWID - 1):0])
    ,.mst5_awlen(mst5_awlen[7:0])
    ,.mst5_awready(mst5_awready)
    ,.mst5_awvalid(mst5_awvalid)
    ,.mst5_bid(mst5_bid[(IDWID - 1):0])
    ,.mst5_bready(mst5_bready)
    ,.mst5_bresp(mst5_bresp[1:0])
    ,.mst5_bvalid(mst5_bvalid)
    ,.mst5_rdata(mst5_rdata[(DWID - 1):0])
    ,.mst5_rid(mst5_rid[(IDWID - 1):0])
    ,.mst5_rlast(mst5_rlast)
    ,.mst5_rready(mst5_rready)
    ,.mst5_rresp(mst5_rresp[1:0])
    ,.mst5_rvalid(mst5_rvalid)
    ,.mst5_wdata(mst5_wdata[(DWID - 1):0])
    ,.mst5_wlast(mst5_wlast)
    ,.mst5_wready(mst5_wready)
    ,.mst5_wstrb(mst5_wstrb[(WSTRB - 1):0])
    ,.mst5_wvalid(mst5_wvalid)

    ,.mst6_araddr(mst6_araddr[31:0])
    ,.mst6_arburst(mst6_arburst[1:0])
    ,.mst6_arextras(mst6_arextras[(EXTRAS - 1):0])
    ,.mst6_arid(mst6_arid[(IDWID - 1):0])
    ,.mst6_arlen(mst6_arlen[7:0])
    ,.mst6_arready(mst6_arready)
    ,.mst6_arvalid(mst6_arvalid)
    ,.mst6_awaddr(mst6_awaddr[31:0])
    ,.mst6_awburst(mst6_awburst[1:0])
    ,.mst6_awextras(mst6_awextras[(EXTRAS - 1):0])
    ,.mst6_awid(mst6_awid[(IDWID - 1):0])
    ,.mst6_awlen(mst6_awlen[7:0])
    ,.mst6_awready(mst6_awready)
    ,.mst6_awvalid(mst6_awvalid)
    ,.mst6_bid(mst6_bid[(IDWID - 1):0])
    ,.mst6_bready(mst6_bready)
    ,.mst6_bresp(mst6_bresp[1:0])
    ,.mst6_bvalid(mst6_bvalid)
    ,.mst6_rdata(mst6_rdata[(DWID - 1):0])
    ,.mst6_rid(mst6_rid[(IDWID - 1):0])
    ,.mst6_rlast(mst6_rlast)
    ,.mst6_rready(mst6_rready)
    ,.mst6_rresp(mst6_rresp[1:0])
    ,.mst6_rvalid(mst6_rvalid)
    ,.mst6_wdata(mst6_wdata[(DWID - 1):0])
    ,.mst6_wlast(mst6_wlast)
    ,.mst6_wready(mst6_wready)
    ,.mst6_wstrb(mst6_wstrb[(WSTRB - 1):0])
    ,.mst6_wvalid(mst6_wvalid)

    ,.mst7_araddr(mst7_araddr[31:0])
    ,.mst7_arburst(mst7_arburst[1:0])
    ,.mst7_arextras(mst7_arextras[(EXTRAS - 1):0])
    ,.mst7_arid(mst7_arid[(IDWID - 1):0])
    ,.mst7_arlen(mst7_arlen[7:0])
    ,.mst7_arready(mst7_arready)
    ,.mst7_arvalid(mst7_arvalid)
    ,.mst7_awaddr(mst7_awaddr[31:0])
    ,.mst7_awburst(mst7_awburst[1:0])
    ,.mst7_awextras(mst7_awextras[(EXTRAS - 1):0])
    ,.mst7_awid(mst7_awid[(IDWID - 1):0])
    ,.mst7_awlen(mst7_awlen[7:0])
    ,.mst7_awready(mst7_awready)
    ,.mst7_awvalid(mst7_awvalid)
    ,.mst7_bid(mst7_bid[(IDWID - 1):0])
    ,.mst7_bready(mst7_bready)
    ,.mst7_bresp(mst7_bresp[1:0])
    ,.mst7_bvalid(mst7_bvalid)
    ,.mst7_rdata(mst7_rdata[(DWID - 1):0])
    ,.mst7_rid(mst7_rid[(IDWID - 1):0])
    ,.mst7_rlast(mst7_rlast)
    ,.mst7_rready(mst7_rready)
    ,.mst7_rresp(mst7_rresp[1:0])
    ,.mst7_rvalid(mst7_rvalid)
    ,.mst7_wdata(mst7_wdata[(DWID - 1):0])
    ,.mst7_wlast(mst7_wlast)
    ,.mst7_wready(mst7_wready)
    ,.mst7_wstrb(mst7_wstrb[(WSTRB - 1):0])
    ,.mst7_wvalid(mst7_wvalid)

    ,.mst8_araddr(mst8_araddr[31:0])
    ,.mst8_arburst(mst8_arburst[1:0])
    ,.mst8_arextras(mst8_arextras[(EXTRAS - 1):0])
    ,.mst8_arid(mst8_arid[(IDWID - 1):0])
    ,.mst8_arlen(mst8_arlen[7:0])
    ,.mst8_arready(mst8_arready)
    ,.mst8_arvalid(mst8_arvalid)
    ,.mst8_awaddr(mst8_awaddr[31:0])
    ,.mst8_awburst(mst8_awburst[1:0])
    ,.mst8_awextras(mst8_awextras[(EXTRAS - 1):0])
    ,.mst8_awid(mst8_awid[(IDWID - 1):0])
    ,.mst8_awlen(mst8_awlen[7:0])
    ,.mst8_awready(mst8_awready)
    ,.mst8_awvalid(mst8_awvalid)
    ,.mst8_bid(mst8_bid[(IDWID - 1):0])
    ,.mst8_bready(mst8_bready)
    ,.mst8_bresp(mst8_bresp[1:0])
    ,.mst8_bvalid(mst8_bvalid)
    ,.mst8_rdata(mst8_rdata[(DWID - 1):0])
    ,.mst8_rid(mst8_rid[(IDWID - 1):0])
    ,.mst8_rlast(mst8_rlast)
    ,.mst8_rready(mst8_rready)
    ,.mst8_rresp(mst8_rresp[1:0])
    ,.mst8_rvalid(mst8_rvalid)
    ,.mst8_wdata(mst8_wdata[(DWID - 1):0])
    ,.mst8_wlast(mst8_wlast)
    ,.mst8_wready(mst8_wready)
    ,.mst8_wstrb(mst8_wstrb[(WSTRB - 1):0])
    ,.mst8_wvalid(mst8_wvalid)

    ,.mst9_araddr(mst9_araddr[31:0])
    ,.mst9_arburst(mst9_arburst[1:0])
    ,.mst9_arextras(mst9_arextras[(EXTRAS - 1):0])
    ,.mst9_arid(mst9_arid[(IDWID - 1):0])
    ,.mst9_arlen(mst9_arlen[7:0])
    ,.mst9_arready(mst9_arready)
    ,.mst9_arvalid(mst9_arvalid)
    ,.mst9_awaddr(mst9_awaddr[31:0])
    ,.mst9_awburst(mst9_awburst[1:0])
    ,.mst9_awextras(mst9_awextras[(EXTRAS - 1):0])
    ,.mst9_awid(mst9_awid[(IDWID - 1):0])
    ,.mst9_awlen(mst9_awlen[7:0])
    ,.mst9_awready(mst9_awready)
    ,.mst9_awvalid(mst9_awvalid)
    ,.mst9_bid(mst9_bid[(IDWID - 1):0])
    ,.mst9_bready(mst9_bready)
    ,.mst9_bresp(mst9_bresp[1:0])
    ,.mst9_bvalid(mst9_bvalid)
    ,.mst9_rdata(mst9_rdata[(DWID - 1):0])
    ,.mst9_rid(mst9_rid[(IDWID - 1):0])
    ,.mst9_rlast(mst9_rlast)
    ,.mst9_rready(mst9_rready)
    ,.mst9_rresp(mst9_rresp[1:0])
    ,.mst9_rvalid(mst9_rvalid)
    ,.mst9_wdata(mst9_wdata[(DWID - 1):0])
    ,.mst9_wlast(mst9_wlast)
    ,.mst9_wready(mst9_wready)
    ,.mst9_wstrb(mst9_wstrb[(WSTRB - 1):0])
    ,.mst9_wvalid(mst9_wvalid)
);
endmodule
