`define NC100_RGF_BASEADDR    'h0
`define ADDR_REGA                                                'h0
`define ADDR_CONTROL0                                            'h4
`define ADDR_STATUSA                                             'h8
`define ADDR_REGB                                                'hc
`define ADDR_EXTERN                                              'h10
`define ADDR_LDST_RAM                                            'h800
