module logtab ( input [9:0] index,output [31:0] result);
assign result = 
    (index==0) ? 32'h00000000 : // 0.0 
    (index==1) ? 32'h3ab89200 : // 0.00140819439281 
    (index==2) ? 32'h3b387c00 : // 0.00281501560705 
    (index==3) ? 32'h3b8a4b80 : // 0.0042204663182 
    (index==4) ? 32'h3bb84e00 : // 0.00562454919388 
    (index==5) ? 32'h3be64480 : // 0.00702726689397 
    (index==6) ? 32'h3c0a1800 : // 0.00842862207058 
    (index==7) ? 32'h3c210800 : // 0.00982861736811 
    (index==8) ? 32'h3c37f280 : // 0.0112272554233 
    (index==9) ? 32'h3c4ed700 : // 0.0126245388651 
    (index==10) ? 32'h3c65b600 : // 0.0140204703149 
    (index==11) ? 32'h3c7c8f40 : // 0.0154150523867 
    (index==12) ? 32'h3c89b180 : // 0.0168082876866 
    (index==13) ? 32'h3c951880 : // 0.0182001788132 
    (index==14) ? 32'h3ca07ca0 : // 0.0195907283579 
    (index==15) ? 32'h3cabde00 : // 0.0209799389042 
    (index==16) ? 32'h3cb73ca0 : // 0.0223678130285 
    (index==17) ? 32'h3cc29860 : // 0.0237543532994 
    (index==18) ? 32'h3ccdf160 : // 0.0251395622785 
    (index==19) ? 32'h3cd947a0 : // 0.0265234425198 
    (index==20) ? 32'h3ce49b00 : // 0.0279059965699 
    (index==21) ? 32'h3cefebc0 : // 0.0292872269682 
    (index==22) ? 32'h3cfb39a0 : // 0.0306671362469 
    (index==23) ? 32'h3d034260 : // 0.0320457269308 
    (index==24) ? 32'h3d08e680 : // 0.0334230015375 
    (index==25) ? 32'h3d0e8950 : // 0.0347989625773 
    (index==26) ? 32'h3d142ac0 : // 0.0361736125535 
    (index==27) ? 32'h3d19cad0 : // 0.0375469539622 
    (index==28) ? 32'h3d1f6980 : // 0.0389189892923 
    (index==29) ? 32'h3d2506d0 : // 0.0402897210257 
    (index==30) ? 32'h3d2aa2c0 : // 0.0416591516372 
    (index==31) ? 32'h3d303d60 : // 0.0430272835945 
    (index==32) ? 32'h3d35d690 : // 0.0443941193585 
    (index==33) ? 32'h3d3b6e70 : // 0.0457596613827 
    (index==34) ? 32'h3d410500 : // 0.047123912114 
    (index==35) ? 32'h3d469a20 : // 0.0484868739923 
    (index==36) ? 32'h3d4c2df0 : // 0.0498485494506 
    (index==37) ? 32'h3d51c070 : // 0.0512089409148 
    (index==38) ? 32'h3d575190 : // 0.0525680508042 
    (index==39) ? 32'h3d5ce160 : // 0.0539258815311 
    (index==40) ? 32'h3d626fd0 : // 0.0552824355012 
    (index==41) ? 32'h3d67fcf0 : // 0.0566377151132 
    (index==42) ? 32'h3d6d88b0 : // 0.0579917227592 
    (index==43) ? 32'h3d731320 : // 0.0593444608244 
    (index==44) ? 32'h3d789c40 : // 0.0606959316876 
    (index==45) ? 32'h3d7e2410 : // 0.0620461377205 
    (index==46) ? 32'h3d81d540 : // 0.0633950812885 
    (index==47) ? 32'h3d8497d8 : // 0.0647427647503 
    (index==48) ? 32'h3d8759c0 : // 0.0660891904578 
    (index==49) ? 32'h3d8a1b00 : // 0.0674343607565 
    (index==50) ? 32'h3d8cdba0 : // 0.0687782779854 
    (index==51) ? 32'h3d8f9b90 : // 0.0701209444768 
    (index==52) ? 32'h3d925ad8 : // 0.0714623625566 
    (index==53) ? 32'h3d951978 : // 0.0728025345442 
    (index==54) ? 32'h3d97d778 : // 0.0741414627525 
    (index==55) ? 32'h3d9a94c8 : // 0.075479149488 
    (index==56) ? 32'h3d9d5178 : // 0.0768155970508 
    (index==57) ? 32'h3da00d80 : // 0.0781508077347 
    (index==58) ? 32'h3da2c8e8 : // 0.0794847838268 
    (index==59) ? 32'h3da583a8 : // 0.0808175276083 
    (index==60) ? 32'h3da83dc0 : // 0.0821490413539 
    (index==61) ? 32'h3daaf730 : // 0.0834793273318 
    (index==62) ? 32'h3dadb000 : // 0.0848083878044 
    (index==63) ? 32'h3db06830 : // 0.0861362250273 
    (index==64) ? 32'h3db31fb0 : // 0.0874628412503 
    (index==65) ? 32'h3db5d698 : // 0.0887882387169 
    (index==66) ? 32'h3db88cd8 : // 0.0901124196643 
    (index==67) ? 32'h3dbb4278 : // 0.0914353863236 
    (index==68) ? 32'h3dbdf770 : // 0.0927571409199 
    (index==69) ? 32'h3dc0abc8 : // 0.0940776856719 
    (index==70) ? 32'h3dc35f80 : // 0.0953970227926 
    (index==71) ? 32'h3dc61298 : // 0.0967151544885 
    (index==72) ? 32'h3dc8c508 : // 0.0980320829605 
    (index==73) ? 32'h3dcb76d8 : // 0.0993478104032 
    (index==74) ? 32'h3dce2808 : // 0.100662339005 
    (index==75) ? 32'h3dd0d898 : // 0.101975670949 
    (index==76) ? 32'h3dd38888 : // 0.103287808412 
    (index==77) ? 32'h3dd637d8 : // 0.104598753564 
    (index==78) ? 32'h3dd8e688 : // 0.105908508571 
    (index==79) ? 32'h3ddb94a0 : // 0.107217075591 
    (index==80) ? 32'h3dde4210 : // 0.108524456778 
    (index==81) ? 32'h3de0eee0 : // 0.109830654279 
    (index==82) ? 32'h3de39b18 : // 0.111135670235 
    (index==83) ? 32'h3de646a8 : // 0.112439506782 
    (index==84) ? 32'h3de8f1a0 : // 0.113742166049 
    (index==85) ? 32'h3deb9c00 : // 0.115043650162 
    (index==86) ? 32'h3dee45b8 : // 0.116343961237 
    (index==87) ? 32'h3df0eed8 : // 0.117643101389 
    (index==88) ? 32'h3df39760 : // 0.118941072724 
    (index==89) ? 32'h3df63f40 : // 0.120237877342 
    (index==90) ? 32'h3df8e690 : // 0.12153351734 
    (index==91) ? 32'h3dfb8d38 : // 0.122827994808 
    (index==92) ? 32'h3dfe3350 : // 0.124121311829 
    (index==93) ? 32'h3e006c60 : // 0.125413470483 
    (index==94) ? 32'h3e01bed0 : // 0.126704472843 
    (index==95) ? 32'h3e0310f0 : // 0.127994320976 
    (index==96) ? 32'h3e0462c4 : // 0.129283016945 
    (index==97) ? 32'h3e05b448 : // 0.130570562805 
    (index==98) ? 32'h3e070580 : // 0.131856960609 
    (index==99) ? 32'h3e08566c : // 0.133142212401 
    (index==100) ? 32'h3e09a70c : // 0.134426320221 
    (index==101) ? 32'h3e0af760 : // 0.135709286104 
    (index==102) ? 32'h3e0c4764 : // 0.13699111208 
    (index==103) ? 32'h3e0d971c : // 0.138271800172 
    (index==104) ? 32'h3e0ee68c : // 0.139551352399 
    (index==105) ? 32'h3e1035ac : // 0.140829770773 
    (index==106) ? 32'h3e118480 : // 0.142107057303 
    (index==107) ? 32'h3e12d30c : // 0.14338321399 
    (index==108) ? 32'h3e142148 : // 0.144658242832 
    (index==109) ? 32'h3e156f3c : // 0.145932145821 
    (index==110) ? 32'h3e16bce0 : // 0.147204924942 
    (index==111) ? 32'h3e180a3c : // 0.148476582178 
    (index==112) ? 32'h3e19574c : // 0.149747119505 
    (index==113) ? 32'h3e1aa414 : // 0.151016538892 
    (index==114) ? 32'h3e1bf08c : // 0.152284842307 
    (index==115) ? 32'h3e1d3cbc : // 0.153552031708 
    (index==116) ? 32'h3e1e88a0 : // 0.154818109052 
    (index==117) ? 32'h3e1fd43c : // 0.156083076289 
    (index==118) ? 32'h3e211f8c : // 0.157346935363 
    (index==119) ? 32'h3e226a90 : // 0.158609688214 
    (index==120) ? 32'h3e23b54c : // 0.159871336778 
    (index==121) ? 32'h3e24ffc0 : // 0.161131882984 
    (index==122) ? 32'h3e2649e8 : // 0.162391328757 
    (index==123) ? 32'h3e2793c4 : // 0.163649676016 
    (index==124) ? 32'h3e28dd5c : // 0.164906926676 
    (index==125) ? 32'h3e2a26a4 : // 0.166163082646 
    (index==126) ? 32'h3e2b6fa8 : // 0.167418145832 
    (index==127) ? 32'h3e2cb860 : // 0.168672118132 
    (index==128) ? 32'h3e2e00d0 : // 0.169925001442 
    (index==129) ? 32'h3e2f48f8 : // 0.171176797652 
    (index==130) ? 32'h3e3090d4 : // 0.172427508645 
    (index==131) ? 32'h3e31d868 : // 0.173677136303 
    (index==132) ? 32'h3e331fb4 : // 0.174925682501 
    (index==133) ? 32'h3e3466b8 : // 0.176173149107 
    (index==134) ? 32'h3e35ad74 : // 0.177419537989 
    (index==135) ? 32'h3e36f3e8 : // 0.178664851006 
    (index==136) ? 32'h3e383a14 : // 0.179909090015 
    (index==137) ? 32'h3e397ff8 : // 0.181152256866 
    (index==138) ? 32'h3e3ac594 : // 0.182394353405 
    (index==139) ? 32'h3e3c0ae8 : // 0.183635381473 
    (index==140) ? 32'h3e3d4ff4 : // 0.184875342908 
    (index==141) ? 32'h3e3e94b8 : // 0.186114239542 
    (index==142) ? 32'h3e3fd938 : // 0.1873520732 
    (index==143) ? 32'h3e411d6c : // 0.188588845707 
    (index==144) ? 32'h3e42615c : // 0.18982455888 
    (index==145) ? 32'h3e43a504 : // 0.191059214532 
    (index==146) ? 32'h3e44e868 : // 0.192292814471 
    (index==147) ? 32'h3e462b80 : // 0.193525360501 
    (index==148) ? 32'h3e476e54 : // 0.194756854422 
    (index==149) ? 32'h3e48b0e4 : // 0.195987298029 
    (index==150) ? 32'h3e49f32c : // 0.19721669311 
    (index==151) ? 32'h3e4b352c : // 0.198445041452 
    (index==152) ? 32'h3e4c76e8 : // 0.199672344836 
    (index==153) ? 32'h3e4db85c : // 0.200898605038 
    (index==154) ? 32'h3e4ef98c : // 0.20212382383 
    (index==155) ? 32'h3e503a74 : // 0.20334800298 
    (index==156) ? 32'h3e517b18 : // 0.204571144249 
    (index==157) ? 32'h3e52bb74 : // 0.205793249397 
    (index==158) ? 32'h3e53fb8c : // 0.207014320178 
    (index==159) ? 32'h3e553b60 : // 0.20823435834 
    (index==160) ? 32'h3e567af0 : // 0.209453365629 
    (index==161) ? 32'h3e57ba38 : // 0.210671343786 
    (index==162) ? 32'h3e58f93c : // 0.211888294546 
    (index==163) ? 32'h3e5a37fc : // 0.213104219642 
    (index==164) ? 32'h3e5b7678 : // 0.214319120801 
    (index==165) ? 32'h3e5cb4ac : // 0.215532999746 
    (index==166) ? 32'h3e5df2a0 : // 0.216745858195 
    (index==167) ? 32'h3e5f304c : // 0.217957697864 
    (index==168) ? 32'h3e606db4 : // 0.219168520462 
    (index==169) ? 32'h3e61aad8 : // 0.220378327695 
    (index==170) ? 32'h3e62e7b8 : // 0.221587121265 
    (index==171) ? 32'h3e642458 : // 0.222794902868 
    (index==172) ? 32'h3e6560b0 : // 0.224001674198 
    (index==173) ? 32'h3e669cc4 : // 0.225207436944 
    (index==174) ? 32'h3e67d898 : // 0.226412192789 
    (index==175) ? 32'h3e691424 : // 0.227615943414 
    (index==176) ? 32'h3e6a4f70 : // 0.228818690496 
    (index==177) ? 32'h3e6b8a78 : // 0.230020435706 
    (index==178) ? 32'h3e6cc53c : // 0.231221180711 
    (index==179) ? 32'h3e6dffc0 : // 0.232420927176 
    (index==180) ? 32'h3e6f39fc : // 0.23361967676 
    (index==181) ? 32'h3e7073f8 : // 0.234817431117 
    (index==182) ? 32'h3e71adb4 : // 0.2360141919 
    (index==183) ? 32'h3e72e728 : // 0.237209960755 
    (index==184) ? 32'h3e74205c : // 0.238404739325 
    (index==185) ? 32'h3e755950 : // 0.239598529249 
    (index==186) ? 32'h3e769200 : // 0.240791332162 
    (index==187) ? 32'h3e77ca6c : // 0.241983149694 
    (index==188) ? 32'h3e790298 : // 0.243173983473 
    (index==189) ? 32'h3e7a3a80 : // 0.244363835121 
    (index==190) ? 32'h3e7b7228 : // 0.245552706256 
    (index==191) ? 32'h3e7ca990 : // 0.246740598493 
    (index==192) ? 32'h3e7de0b4 : // 0.247927513444 
    (index==193) ? 32'h3e7f1798 : // 0.249113452714 
    (index==194) ? 32'h3e80271c : // 0.250298417906 
    (index==195) ? 32'h3e80c24c : // 0.25148241062 
    (index==196) ? 32'h3e815d5c : // 0.25266543245 
    (index==197) ? 32'h3e81f84c : // 0.253847484987 
    (index==198) ? 32'h3e82931a : // 0.255028569819 
    (index==199) ? 32'h3e832dc8 : // 0.256208688527 
    (index==200) ? 32'h3e83c856 : // 0.257387842693 
    (index==201) ? 32'h3e8462c4 : // 0.25856603389 
    (index==202) ? 32'h3e84fd10 : // 0.259743263691 
    (index==203) ? 32'h3e85973e : // 0.260919533663 
    (index==204) ? 32'h3e86314a : // 0.26209484537 
    (index==205) ? 32'h3e86cb38 : // 0.263269200373 
    (index==206) ? 32'h3e876504 : // 0.264442600227 
    (index==207) ? 32'h3e87feb2 : // 0.265615046484 
    (index==208) ? 32'h3e88983e : // 0.266786540695 
    (index==209) ? 32'h3e8931aa : // 0.267957084403 
    (index==210) ? 32'h3e89caf8 : // 0.269126679149 
    (index==211) ? 32'h3e8a6426 : // 0.270295326472 
    (index==212) ? 32'h3e8afd32 : // 0.271463027904 
    (index==213) ? 32'h3e8b9620 : // 0.272629784976 
    (index==214) ? 32'h3e8c2eee : // 0.273795599214 
    (index==215) ? 32'h3e8cc79e : // 0.274960472141 
    (index==216) ? 32'h3e8d602c : // 0.276124405274 
    (index==217) ? 32'h3e8df89c : // 0.27728740013 
    (index==218) ? 32'h3e8e90ec : // 0.27844945822 
    (index==219) ? 32'h3e8f291e : // 0.279610581052 
    (index==220) ? 32'h3e8fc12e : // 0.280770770131 
    (index==221) ? 32'h3e905920 : // 0.281930026955 
    (index==222) ? 32'h3e90f0f4 : // 0.283088353024 
    (index==223) ? 32'h3e9188a8 : // 0.28424574983 
    (index==224) ? 32'h3e92203c : // 0.285402218862 
    (index==225) ? 32'h3e92b7b2 : // 0.286557761608 
    (index==226) ? 32'h3e934f08 : // 0.287712379549 
    (index==227) ? 32'h3e93e640 : // 0.288866074166 
    (index==228) ? 32'h3e947d58 : // 0.290018846933 
    (index==229) ? 32'h3e951452 : // 0.291170699322 
    (index==230) ? 32'h3e95ab2e : // 0.292321632802 
    (index==231) ? 32'h3e9641ea : // 0.293471648838 
    (index==232) ? 32'h3e96d886 : // 0.294620748892 
    (index==233) ? 32'h3e976f06 : // 0.295768934421 
    (index==234) ? 32'h3e980566 : // 0.296916206879 
    (index==235) ? 32'h3e989ba8 : // 0.298062567719 
    (index==236) ? 32'h3e9931ca : // 0.299208018387 
    (index==237) ? 32'h3e99c7ce : // 0.300352560328 
    (index==238) ? 32'h3e9a5db4 : // 0.301496194983 
    (index==239) ? 32'h3e9af37c : // 0.302638923788 
    (index==240) ? 32'h3e9b8926 : // 0.303780748177 
    (index==241) ? 32'h3e9c1eb0 : // 0.304921669582 
    (index==242) ? 32'h3e9cb41e : // 0.306061689428 
    (index==243) ? 32'h3e9d496c : // 0.307200809141 
    (index==244) ? 32'h3e9dde9c : // 0.308339030139 
    (index==245) ? 32'h3e9e73ae : // 0.309476353841 
    (index==246) ? 32'h3e9f08a2 : // 0.31061278166 
    (index==247) ? 32'h3e9f9d78 : // 0.311748315005 
    (index==248) ? 32'h3ea03230 : // 0.312882955284 
    (index==249) ? 32'h3ea0c6cc : // 0.314016703901 
    (index==250) ? 32'h3ea15b48 : // 0.315149562256 
    (index==251) ? 32'h3ea1efa6 : // 0.316281531746 
    (index==252) ? 32'h3ea283e6 : // 0.317412613765 
    (index==253) ? 32'h3ea3180a : // 0.318542809703 
    (index==254) ? 32'h3ea3ac10 : // 0.319672120947 
    (index==255) ? 32'h3ea43ff8 : // 0.320800548882 
    (index==256) ? 32'h3ea4d3c2 : // 0.321928094887 
    (index==257) ? 32'h3ea5676e : // 0.323054760342 
    (index==258) ? 32'h3ea5fafe : // 0.324180546619 
    (index==259) ? 32'h3ea68e6e : // 0.32530545509 
    (index==260) ? 32'h3ea721c4 : // 0.326429487122 
    (index==261) ? 32'h3ea7b4fa : // 0.327552644081 
    (index==262) ? 32'h3ea84814 : // 0.328674927328 
    (index==263) ? 32'h3ea8db10 : // 0.329796338221 
    (index==264) ? 32'h3ea96dee : // 0.330916878115 
    (index==265) ? 32'h3eaa00b0 : // 0.332036548362 
    (index==266) ? 32'h3eaa9356 : // 0.333155350311 
    (index==267) ? 32'h3eab25de : // 0.334273285307 
    (index==268) ? 32'h3eabb848 : // 0.335390354694 
    (index==269) ? 32'h3eac4a96 : // 0.33650655981 
    (index==270) ? 32'h3eacdcc6 : // 0.337621901993 
    (index==271) ? 32'h3ead6eda : // 0.338736382574 
    (index==272) ? 32'h3eae00d0 : // 0.339850002885 
    (index==273) ? 32'h3eae92aa : // 0.340962764252 
    (index==274) ? 32'h3eaf2468 : // 0.342074667999 
    (index==275) ? 32'h3eafb608 : // 0.343185715448 
    (index==276) ? 32'h3eb0478c : // 0.344295907916 
    (index==277) ? 32'h3eb0d8f4 : // 0.345405246718 
    (index==278) ? 32'h3eb16a3e : // 0.346513733166 
    (index==279) ? 32'h3eb1fb6c : // 0.347621368568 
    (index==280) ? 32'h3eb28c7e : // 0.348728154231 
    (index==281) ? 32'h3eb31d74 : // 0.349834091457 
    (index==282) ? 32'h3eb3ae4c : // 0.350939181546 
    (index==283) ? 32'h3eb43f08 : // 0.352043425795 
    (index==284) ? 32'h3eb4cfa8 : // 0.353146825498 
    (index==285) ? 32'h3eb5602c : // 0.354249381945 
    (index==286) ? 32'h3eb5f094 : // 0.355351096425 
    (index==287) ? 32'h3eb680de : // 0.356451970222 
    (index==288) ? 32'h3eb7110e : // 0.357552004618 
    (index==289) ? 32'h3eb7a120 : // 0.358651200893 
    (index==290) ? 32'h3eb83118 : // 0.359749560322 
    (index==291) ? 32'h3eb8c0f2 : // 0.36084708418 
    (index==292) ? 32'h3eb950b0 : // 0.361943773735 
    (index==293) ? 32'h3eb9e054 : // 0.363039630257 
    (index==294) ? 32'h3eba6fda : // 0.364134655008 
    (index==295) ? 32'h3ebaff46 : // 0.365228849252 
    (index==296) ? 32'h3ebb8e94 : // 0.366322214246 
    (index==297) ? 32'h3ebc1dc8 : // 0.367414751247 
    (index==298) ? 32'h3ebcace0 : // 0.368506461508 
    (index==299) ? 32'h3ebd3bdc : // 0.369597346279 
    (index==300) ? 32'h3ebdcabc : // 0.370687406807 
    (index==301) ? 32'h3ebe5982 : // 0.371776644338 
    (index==302) ? 32'h3ebee82a : // 0.372865060113 
    (index==303) ? 32'h3ebf76b8 : // 0.37395265537 
    (index==304) ? 32'h3ec0052a : // 0.375039431347 
    (index==305) ? 32'h3ec09380 : // 0.376125389276 
    (index==306) ? 32'h3ec121bc : // 0.377210530389 
    (index==307) ? 32'h3ec1afdc : // 0.378294855912 
    (index==308) ? 32'h3ec23de0 : // 0.379378367071 
    (index==309) ? 32'h3ec2cbca : // 0.380461065089 
    (index==310) ? 32'h3ec35998 : // 0.381542951185 
    (index==311) ? 32'h3ec3e74a : // 0.382624026575 
    (index==312) ? 32'h3ec474e2 : // 0.383704292474 
    (index==313) ? 32'h3ec50260 : // 0.384783750093 
    (index==314) ? 32'h3ec58fc0 : // 0.385862400641 
    (index==315) ? 32'h3ec61d08 : // 0.386940245324 
    (index==316) ? 32'h3ec6aa32 : // 0.388017285345 
    (index==317) ? 32'h3ec73744 : // 0.389093521904 
    (index==318) ? 32'h3ec7c438 : // 0.3901689562 
    (index==319) ? 32'h3ec85114 : // 0.391243589427 
    (index==320) ? 32'h3ec8ddd4 : // 0.392317422779 
    (index==321) ? 32'h3ec96a78 : // 0.393390457444 
    (index==322) ? 32'h3ec9f702 : // 0.39446269461 
    (index==323) ? 32'h3eca8372 : // 0.395534135462 
    (index==324) ? 32'h3ecb0fc8 : // 0.396604781182 
    (index==325) ? 32'h3ecb9c02 : // 0.397674632948 
    (index==326) ? 32'h3ecc2822 : // 0.398743691938 
    (index==327) ? 32'h3eccb426 : // 0.399811959326 
    (index==328) ? 32'h3ecd4010 : // 0.400879436282 
    (index==329) ? 32'h3ecdcbe0 : // 0.401946123977 
    (index==330) ? 32'h3ece5796 : // 0.403012023575 
    (index==331) ? 32'h3ecee332 : // 0.404077136241 
    (index==332) ? 32'h3ecf6eb2 : // 0.405141463136 
    (index==333) ? 32'h3ecffa1a : // 0.406205005419 
    (index==334) ? 32'h3ed08566 : // 0.407267764245 
    (index==335) ? 32'h3ed11098 : // 0.408329740767 
    (index==336) ? 32'h3ed19bb0 : // 0.409390936138 
    (index==337) ? 32'h3ed226ac : // 0.410451351504 
    (index==338) ? 32'h3ed2b190 : // 0.411510988012 
    (index==339) ? 32'h3ed33c5a : // 0.412569846805 
    (index==340) ? 32'h3ed3c70a : // 0.413627929024 
    (index==341) ? 32'h3ed4519e : // 0.414685235807 
    (index==342) ? 32'h3ed4dc1a : // 0.41574176829 
    (index==343) ? 32'h3ed5667c : // 0.416797527606 
    (index==344) ? 32'h3ed5f0c2 : // 0.417852514886 
    (index==345) ? 32'h3ed67af0 : // 0.418906731258 
    (index==346) ? 32'h3ed70504 : // 0.419960177848 
    (index==347) ? 32'h3ed78efe : // 0.421012855779 
    (index==348) ? 32'h3ed818de : // 0.422064766173 
    (index==349) ? 32'h3ed8a2a6 : // 0.423115910147 
    (index==350) ? 32'h3ed92c52 : // 0.424166288818 
    (index==351) ? 32'h3ed9b5e6 : // 0.425215903299 
    (index==352) ? 32'h3eda3f5e : // 0.426264754702 
    (index==353) ? 32'h3edac8be : // 0.427312844135 
    (index==354) ? 32'h3edb5206 : // 0.428360172704 
    (index==355) ? 32'h3edbdb32 : // 0.429406741514 
    (index==356) ? 32'h3edc6446 : // 0.430452551666 
    (index==357) ? 32'h3edced40 : // 0.431497604258 
    (index==358) ? 32'h3edd7620 : // 0.432541900388 
    (index==359) ? 32'h3eddfee8 : // 0.43358544115 
    (index==360) ? 32'h3ede8796 : // 0.434628227637 
    (index==361) ? 32'h3edf102c : // 0.435670260937 
    (index==362) ? 32'h3edf98a6 : // 0.436711542137 
    (index==363) ? 32'h3ee0210a : // 0.437752072324 
    (index==364) ? 32'h3ee0a952 : // 0.438791852578 
    (index==365) ? 32'h3ee13182 : // 0.439830883981 
    (index==366) ? 32'h3ee1b99a : // 0.440869167611 
    (index==367) ? 32'h3ee24198 : // 0.441906704542 
    (index==368) ? 32'h3ee2c97c : // 0.442943495849 
    (index==369) ? 32'h3ee35148 : // 0.443979542601 
    (index==370) ? 32'h3ee3d8fc : // 0.445014845868 
    (index==371) ? 32'h3ee46096 : // 0.446049406717 
    (index==372) ? 32'h3ee4e816 : // 0.44708322621 
    (index==373) ? 32'h3ee56f80 : // 0.448116305409 
    (index==374) ? 32'h3ee5f6ce : // 0.449148645375 
    (index==375) ? 32'h3ee67e06 : // 0.450180247165 
    (index==376) ? 32'h3ee70524 : // 0.451211111832 
    (index==377) ? 32'h3ee78c28 : // 0.452241240431 
    (index==378) ? 32'h3ee81316 : // 0.453270634011 
    (index==379) ? 32'h3ee899ea : // 0.45429929362 
    (index==380) ? 32'h3ee920a6 : // 0.455327220305 
    (index==381) ? 32'h3ee9a748 : // 0.456354415108 
    (index==382) ? 32'h3eea2dd2 : // 0.457380879073 
    (index==383) ? 32'h3eeab444 : // 0.458406613237 
    (index==384) ? 32'h3eeb3a9e : // 0.459431618637 
    (index==385) ? 32'h3eebc0e0 : // 0.46045589631 
    (index==386) ? 32'h3eec4708 : // 0.461479447286 
    (index==387) ? 32'h3eeccd18 : // 0.462502272597 
    (index==388) ? 32'h3eed5310 : // 0.463524373271 
    (index==389) ? 32'h3eedd8f0 : // 0.464545750334 
    (index==390) ? 32'h3eee5eb8 : // 0.465566404809 
    (index==391) ? 32'h3eeee466 : // 0.466586337719 
    (index==392) ? 32'h3eef69fe : // 0.467605550083 
    (index==393) ? 32'h3eefef7c : // 0.468624042918 
    (index==394) ? 32'h3ef074e4 : // 0.46964181724 
    (index==395) ? 32'h3ef0fa32 : // 0.470658874061 
    (index==396) ? 32'h3ef17f68 : // 0.471675214392 
    (index==397) ? 32'h3ef20488 : // 0.472690839243 
    (index==398) ? 32'h3ef2898e : // 0.473705749619 
    (index==399) ? 32'h3ef30e7e : // 0.474719946526 
    (index==400) ? 32'h3ef39354 : // 0.475733430966 
    (index==401) ? 32'h3ef41814 : // 0.476746203939 
    (index==402) ? 32'h3ef49cba : // 0.477758266444 
    (index==403) ? 32'h3ef5214a : // 0.478769619476 
    (index==404) ? 32'h3ef5a5c2 : // 0.479780264029 
    (index==405) ? 32'h3ef62a22 : // 0.480790201096 
    (index==406) ? 32'h3ef6ae6a : // 0.481799431666 
    (index==407) ? 32'h3ef7329a : // 0.482807956727 
    (index==408) ? 32'h3ef7b6b2 : // 0.483815777264 
    (index==409) ? 32'h3ef83ab4 : // 0.484822894262 
    (index==410) ? 32'h3ef8be9e : // 0.485829308702 
    (index==411) ? 32'h3ef94270 : // 0.486835021563 
    (index==412) ? 32'h3ef9c62a : // 0.487840033823 
    (index==413) ? 32'h3efa49ce : // 0.488844346457 
    (index==414) ? 32'h3efacd5a : // 0.489847960439 
    (index==415) ? 32'h3efb50ce : // 0.49085087674 
    (index==416) ? 32'h3efbd42a : // 0.49185309633 
    (index==417) ? 32'h3efc5770 : // 0.492854620175 
    (index==418) ? 32'h3efcda9e : // 0.493855449241 
    (index==419) ? 32'h3efd5db6 : // 0.494855584491 
    (index==420) ? 32'h3efde0b4 : // 0.495855026887 
    (index==421) ? 32'h3efe639e : // 0.496853777388 
    (index==422) ? 32'h3efee66e : // 0.497851836951 
    (index==423) ? 32'h3eff6928 : // 0.498849206532 
    (index==424) ? 32'h3effebcc : // 0.499845887083 
    (index==425) ? 32'h3f00372c : // 0.500841879557 
    (index==426) ? 32'h3f007866 : // 0.501837184902 
    (index==427) ? 32'h3f00b995 : // 0.502831804067 
    (index==428) ? 32'h3f00fab9 : // 0.503825737996 
    (index==429) ? 32'h3f013bd1 : // 0.504818987633 
    (index==430) ? 32'h3f017cdd : // 0.50581155392 
    (index==431) ? 32'h3f01bdde : // 0.506803437796 
    (index==432) ? 32'h3f01fed4 : // 0.507794640199 
    (index==433) ? 32'h3f023fbe : // 0.508785162065 
    (index==434) ? 32'h3f02809d : // 0.509775004327 
    (index==435) ? 32'h3f02c170 : // 0.510764167918 
    (index==436) ? 32'h3f030238 : // 0.511752653767 
    (index==437) ? 32'h3f0342f5 : // 0.512740462803 
    (index==438) ? 32'h3f0383a6 : // 0.513727595952 
    (index==439) ? 32'h3f03c44c : // 0.514714054138 
    (index==440) ? 32'h3f0404e7 : // 0.515699838284 
    (index==441) ? 32'h3f044576 : // 0.51668494931 
    (index==442) ? 32'h3f0485fb : // 0.517669388134 
    (index==443) ? 32'h3f04c674 : // 0.518653155673 
    (index==444) ? 32'h3f0506e1 : // 0.519636252843 
    (index==445) ? 32'h3f054744 : // 0.520618680556 
    (index==446) ? 32'h3f05879b : // 0.521600439724 
    (index==447) ? 32'h3f05c7e7 : // 0.522581531255 
    (index==448) ? 32'h3f060828 : // 0.523561956057 
    (index==449) ? 32'h3f06485d : // 0.524541715036 
    (index==450) ? 32'h3f068888 : // 0.525520809095 
    (index==451) ? 32'h3f06c8a7 : // 0.526499239137 
    (index==452) ? 32'h3f0708bb : // 0.52747700606 
    (index==453) ? 32'h3f0748c4 : // 0.528454110765 
    (index==454) ? 32'h3f0788c2 : // 0.529430554146 
    (index==455) ? 32'h3f07c8b5 : // 0.530406337099 
    (index==456) ? 32'h3f08089d : // 0.531381460516 
    (index==457) ? 32'h3f08487a : // 0.532355925289 
    (index==458) ? 32'h3f08884c : // 0.533329732306 
    (index==459) ? 32'h3f08c812 : // 0.534302882455 
    (index==460) ? 32'h3f0907ce : // 0.535275376621 
    (index==461) ? 32'h3f09477f : // 0.536247215688 
    (index==462) ? 32'h3f098725 : // 0.537218400539 
    (index==463) ? 32'h3f09c6bf : // 0.538188932052 
    (index==464) ? 32'h3f0a064f : // 0.539158811108 
    (index==465) ? 32'h3f0a45d4 : // 0.540128038582 
    (index==466) ? 32'h3f0a854e : // 0.54109661535 
    (index==467) ? 32'h3f0ac4bd : // 0.542064542283 
    (index==468) ? 32'h3f0b0422 : // 0.543031820255 
    (index==469) ? 32'h3f0b437b : // 0.543998450135 
    (index==470) ? 32'h3f0b82ca : // 0.544964432789 
    (index==471) ? 32'h3f0bc20d : // 0.545929769085 
    (index==472) ? 32'h3f0c0146 : // 0.546894459888 
    (index==473) ? 32'h3f0c4074 : // 0.547858506058 
    (index==474) ? 32'h3f0c7f97 : // 0.548821908459 
    (index==475) ? 32'h3f0cbeb0 : // 0.549784667948 
    (index==476) ? 32'h3f0cfdbd : // 0.550746785383 
    (index==477) ? 32'h3f0d3cc0 : // 0.551708261621 
    (index==478) ? 32'h3f0d7bb8 : // 0.552669097514 
    (index==479) ? 32'h3f0dbaa6 : // 0.553629293916 
    (index==480) ? 32'h3f0df988 : // 0.554588851678 
    (index==481) ? 32'h3f0e3860 : // 0.555547771647 
    (index==482) ? 32'h3f0e772e : // 0.556506054672 
    (index==483) ? 32'h3f0eb5f0 : // 0.557463701598 
    (index==484) ? 32'h3f0ef4a8 : // 0.558420713269 
    (index==485) ? 32'h3f0f3356 : // 0.559377090527 
    (index==486) ? 32'h3f0f71f8 : // 0.560332834212 
    (index==487) ? 32'h3f0fb091 : // 0.561287945165 
    (index==488) ? 32'h3f0fef1e : // 0.562242424221 
    (index==489) ? 32'h3f102da1 : // 0.563196272217 
    (index==490) ? 32'h3f106c19 : // 0.564149489986 
    (index==491) ? 32'h3f10aa87 : // 0.56510207836 
    (index==492) ? 32'h3f10e8ea : // 0.566054038171 
    (index==493) ? 32'h3f112743 : // 0.567005370247 
    (index==494) ? 32'h3f116591 : // 0.567956075415 
    (index==495) ? 32'h3f11a3d5 : // 0.568906154502 
    (index==496) ? 32'h3f11e20e : // 0.569855608331 
    (index==497) ? 32'h3f12203d : // 0.570804437724 
    (index==498) ? 32'h3f125e61 : // 0.571752643504 
    (index==499) ? 32'h3f129c7b : // 0.572700226487 
    (index==500) ? 32'h3f12da8a : // 0.573647187493 
    (index==501) ? 32'h3f13188f : // 0.574593527338 
    (index==502) ? 32'h3f13568a : // 0.575539246835 
    (index==503) ? 32'h3f13947a : // 0.576484346797 
    (index==504) ? 32'h3f13d260 : // 0.577428828036 
    (index==505) ? 32'h3f14103b : // 0.578372691361 
    (index==506) ? 32'h3f144e0c : // 0.57931593758 
    (index==507) ? 32'h3f148bd3 : // 0.5802585675 
    (index==508) ? 32'h3f14c98f : // 0.581200581925 
    (index==509) ? 32'h3f150741 : // 0.582141981659 
    (index==510) ? 32'h3f1544e9 : // 0.583082767503 
    (index==511) ? 32'h3f158287 : // 0.584022940258 
    (index==512) ? 32'h3f15c01a : // 0.584962500721 
    (index==513) ? 32'h3f15fda3 : // 0.585901449691 
    (index==514) ? 32'h3f163b21 : // 0.586839787962 
    (index==515) ? 32'h3f167896 : // 0.587777516328 
    (index==516) ? 32'h3f16b600 : // 0.588714635582 
    (index==517) ? 32'h3f16f360 : // 0.589651146515 
    (index==518) ? 32'h3f1730b6 : // 0.590587049915 
    (index==519) ? 32'h3f176e02 : // 0.591522346571 
    (index==520) ? 32'h3f17ab43 : // 0.592457037268 
    (index==521) ? 32'h3f17e87b : // 0.593391122792 
    (index==522) ? 32'h3f1825a8 : // 0.594324603925 
    (index==523) ? 32'h3f1862cb : // 0.595257481449 
    (index==524) ? 32'h3f189fe4 : // 0.596189756144 
    (index==525) ? 32'h3f18dcf3 : // 0.59712142879 
    (index==526) ? 32'h3f1919f7 : // 0.598052500162 
    (index==527) ? 32'h3f1956f2 : // 0.598982971036 
    (index==528) ? 32'h3f1993e3 : // 0.599912842187 
    (index==529) ? 32'h3f19d0c9 : // 0.600842114387 
    (index==530) ? 32'h3f1a0da6 : // 0.601770788408 
    (index==531) ? 32'h3f1a4a79 : // 0.602698865018 
    (index==532) ? 32'h3f1a8741 : // 0.603626344986 
    (index==533) ? 32'h3f1ac400 : // 0.604553229079 
    (index==534) ? 32'h3f1b00b4 : // 0.605479518062 
    (index==535) ? 32'h3f1b3d5f : // 0.606405212698 
    (index==536) ? 32'h3f1b79ff : // 0.60733031375 
    (index==537) ? 32'h3f1bb696 : // 0.608254821978 
    (index==538) ? 32'h3f1bf323 : // 0.609178738142 
    (index==539) ? 32'h3f1c2fa6 : // 0.610102063 
    (index==540) ? 32'h3f1c6c1f : // 0.611024797307 
    (index==541) ? 32'h3f1ca88e : // 0.61194694182 
    (index==542) ? 32'h3f1ce4f3 : // 0.612868497291 
    (index==543) ? 32'h3f1d214e : // 0.613789464473 
    (index==544) ? 32'h3f1d5d9f : // 0.614709844115 
    (index==545) ? 32'h3f1d99e7 : // 0.615629636968 
    (index==546) ? 32'h3f1dd625 : // 0.616548843779 
    (index==547) ? 32'h3f1e1259 : // 0.617467465294 
    (index==548) ? 32'h3f1e4e83 : // 0.618385502259 
    (index==549) ? 32'h3f1e8aa3 : // 0.619302955416 
    (index==550) ? 32'h3f1ec6b9 : // 0.620219825507 
    (index==551) ? 32'h3f1f02c6 : // 0.621136113275 
    (index==552) ? 32'h3f1f3ec9 : // 0.622051819456 
    (index==553) ? 32'h3f1f7ac2 : // 0.622966944791 
    (index==554) ? 32'h3f1fb6b2 : // 0.623881490013 
    (index==555) ? 32'h3f1ff298 : // 0.62479545586 
    (index==556) ? 32'h3f202e74 : // 0.625708843064 
    (index==557) ? 32'h3f206a46 : // 0.626621652358 
    (index==558) ? 32'h3f20a60f : // 0.627533884473 
    (index==559) ? 32'h3f20e1ce : // 0.628445540137 
    (index==560) ? 32'h3f211d83 : // 0.62935662008 
    (index==561) ? 32'h3f21592f : // 0.630267125027 
    (index==562) ? 32'h3f2194d1 : // 0.631177055704 
    (index==563) ? 32'h3f21d06a : // 0.632086412835 
    (index==564) ? 32'h3f220bf9 : // 0.632995197143 
    (index==565) ? 32'h3f22477e : // 0.633903409349 
    (index==566) ? 32'h3f2282fa : // 0.634811050172 
    (index==567) ? 32'h3f22be6c : // 0.635718120331 
    (index==568) ? 32'h3f22f9d4 : // 0.636624620544 
    (index==569) ? 32'h3f233533 : // 0.637530551525 
    (index==570) ? 32'h3f237089 : // 0.63843591399 
    (index==571) ? 32'h3f23abd5 : // 0.639340708652 
    (index==572) ? 32'h3f23e717 : // 0.640244936222 
    (index==573) ? 32'h3f242250 : // 0.641148597411 
    (index==574) ? 32'h3f245d7f : // 0.642051692928 
    (index==575) ? 32'h3f2498a5 : // 0.64295422348 
    (index==576) ? 32'h3f24d3c2 : // 0.643856189775 
    (index==577) ? 32'h3f250ed5 : // 0.644757592516 
    (index==578) ? 32'h3f2549de : // 0.645658432409 
    (index==579) ? 32'h3f2584df : // 0.646558710155 
    (index==580) ? 32'h3f25bfd5 : // 0.647458426455 
    (index==581) ? 32'h3f25fac3 : // 0.64835758201 
    (index==582) ? 32'h3f2635a7 : // 0.649256177517 
    (index==583) ? 32'h3f267081 : // 0.650154213675 
    (index==584) ? 32'h3f26ab52 : // 0.651051691179 
    (index==585) ? 32'h3f26e61a : // 0.651948610723 
    (index==586) ? 32'h3f2720d9 : // 0.652844973002 
    (index==587) ? 32'h3f275b8e : // 0.653740778707 
    (index==588) ? 32'h3f27963a : // 0.654636028528 
    (index==589) ? 32'h3f27d0dc : // 0.655530723156 
    (index==590) ? 32'h3f280b75 : // 0.656424863278 
    (index==591) ? 32'h3f284605 : // 0.657318449581 
    (index==592) ? 32'h3f28808c : // 0.658211482752 
    (index==593) ? 32'h3f28bb09 : // 0.659103963474 
    (index==594) ? 32'h3f28f57d : // 0.65999589243 
    (index==595) ? 32'h3f292fe8 : // 0.660887270303 
    (index==596) ? 32'h3f296a4a : // 0.661778097772 
    (index==597) ? 32'h3f29a4a2 : // 0.662668375518 
    (index==598) ? 32'h3f29def1 : // 0.663558104217 
    (index==599) ? 32'h3f2a1937 : // 0.664447284548 
    (index==600) ? 32'h3f2a5374 : // 0.665335917185 
    (index==601) ? 32'h3f2a8da7 : // 0.666224002803 
    (index==602) ? 32'h3f2ac7d2 : // 0.667111542075 
    (index==603) ? 32'h3f2b01f3 : // 0.667998535673 
    (index==604) ? 32'h3f2b3c0b : // 0.668884984266 
    (index==605) ? 32'h3f2b761a : // 0.669770888526 
    (index==606) ? 32'h3f2bb020 : // 0.670656249118 
    (index==607) ? 32'h3f2bea1d : // 0.671541066712 
    (index==608) ? 32'h3f2c2411 : // 0.672425341971 
    (index==609) ? 32'h3f2c5dfb : // 0.673309075562 
    (index==610) ? 32'h3f2c97dd : // 0.674192268146 
    (index==611) ? 32'h3f2cd1b5 : // 0.675074920385 
    (index==612) ? 32'h3f2d0b85 : // 0.675957032942 
    (index==613) ? 32'h3f2d454b : // 0.676838606474 
    (index==614) ? 32'h3f2d7f08 : // 0.677719641641 
    (index==615) ? 32'h3f2db8bd : // 0.678600139099 
    (index==616) ? 32'h3f2df268 : // 0.679480099505 
    (index==617) ? 32'h3f2e2c0a : // 0.680359523514 
    (index==618) ? 32'h3f2e65a3 : // 0.681238411778 
    (index==619) ? 32'h3f2e9f34 : // 0.68211676495 
    (index==620) ? 32'h3f2ed8bb : // 0.682994583682 
    (index==621) ? 32'h3f2f123a : // 0.683871868623 
    (index==622) ? 32'h3f2f4baf : // 0.684748620422 
    (index==623) ? 32'h3f2f851c : // 0.685624839726 
    (index==624) ? 32'h3f2fbe7f : // 0.686500527183 
    (index==625) ? 32'h3f2ff7da : // 0.687375683437 
    (index==626) ? 32'h3f30312c : // 0.688250309133 
    (index==627) ? 32'h3f306a74 : // 0.689124404913 
    (index==628) ? 32'h3f30a3b5 : // 0.689997971419 
    (index==629) ? 32'h3f30dcec : // 0.690871009292 
    (index==630) ? 32'h3f31161a : // 0.691743519171 
    (index==631) ? 32'h3f314f3f : // 0.692615501695 
    (index==632) ? 32'h3f31885c : // 0.693486957499 
    (index==633) ? 32'h3f31c170 : // 0.694357887221 
    (index==634) ? 32'h3f31fa7b : // 0.695228291496 
    (index==635) ? 32'h3f32337d : // 0.696098170956 
    (index==636) ? 32'h3f326c76 : // 0.696967526234 
    (index==637) ? 32'h3f32a567 : // 0.697836357962 
    (index==638) ? 32'h3f32de4f : // 0.69870466677 
    (index==639) ? 32'h3f33172e : // 0.699572453287 
    (index==640) ? 32'h3f335004 : // 0.700439718141 
    (index==641) ? 32'h3f3388d1 : // 0.701306461959 
    (index==642) ? 32'h3f33c196 : // 0.702172685366 
    (index==643) ? 32'h3f33fa52 : // 0.703038388986 
    (index==644) ? 32'h3f343306 : // 0.703903573445 
    (index==645) ? 32'h3f346bb0 : // 0.704768239363 
    (index==646) ? 32'h3f34a452 : // 0.705632387361 
    (index==647) ? 32'h3f34dcec : // 0.706496018061 
    (index==648) ? 32'h3f35157c : // 0.707359132081 
    (index==649) ? 32'h3f354e04 : // 0.708221730038 
    (index==650) ? 32'h3f358684 : // 0.70908381255 
    (index==651) ? 32'h3f35befa : // 0.709945380232 
    (index==652) ? 32'h3f35f769 : // 0.710806433699 
    (index==653) ? 32'h3f362fce : // 0.711666973564 
    (index==654) ? 32'h3f36682b : // 0.71252700044 
    (index==655) ? 32'h3f36a07f : // 0.713386514937 
    (index==656) ? 32'h3f36d8cb : // 0.714245517666 
    (index==657) ? 32'h3f37110e : // 0.715104009236 
    (index==658) ? 32'h3f374948 : // 0.715961990255 
    (index==659) ? 32'h3f37817a : // 0.71681946133 
    (index==660) ? 32'h3f37b9a4 : // 0.717676423066 
    (index==661) ? 32'h3f37f1c5 : // 0.718532876069 
    (index==662) ? 32'h3f3829dd : // 0.719388820942 
    (index==663) ? 32'h3f3861ed : // 0.720244258288 
    (index==664) ? 32'h3f3899f4 : // 0.721099188707 
    (index==665) ? 32'h3f38d1f3 : // 0.721953612801 
    (index==666) ? 32'h3f3909ea : // 0.72280753117 
    (index==667) ? 32'h3f3941d7 : // 0.72366094441 
    (index==668) ? 32'h3f3979bd : // 0.72451385312 
    (index==669) ? 32'h3f39b19a : // 0.725366257896 
    (index==670) ? 32'h3f39e96e : // 0.726218159332 
    (index==671) ? 32'h3f3a213b : // 0.727069558024 
    (index==672) ? 32'h3f3a58fe : // 0.727920454563 
    (index==673) ? 32'h3f3a90b9 : // 0.728770849543 
    (index==674) ? 32'h3f3ac86c : // 0.729620743553 
    (index==675) ? 32'h3f3b0017 : // 0.730470137184 
    (index==676) ? 32'h3f3b37b9 : // 0.731319031025 
    (index==677) ? 32'h3f3b6f53 : // 0.732167425663 
    (index==678) ? 32'h3f3ba6e4 : // 0.733015321686 
    (index==679) ? 32'h3f3bde6d : // 0.733862719679 
    (index==680) ? 32'h3f3c15ed : // 0.734709620226 
    (index==681) ? 32'h3f3c4d66 : // 0.735556023912 
    (index==682) ? 32'h3f3c84d6 : // 0.736401931318 
    (index==683) ? 32'h3f3cbc3d : // 0.737247343028 
    (index==684) ? 32'h3f3cf39d : // 0.73809225962 
    (index==685) ? 32'h3f3d2af4 : // 0.738936681676 
    (index==686) ? 32'h3f3d6243 : // 0.739780609773 
    (index==687) ? 32'h3f3d9989 : // 0.740624044489 
    (index==688) ? 32'h3f3dd0c7 : // 0.741466986401 
    (index==689) ? 32'h3f3e07fd : // 0.742309436084 
    (index==690) ? 32'h3f3e3f2b : // 0.743151394112 
    (index==691) ? 32'h3f3e7650 : // 0.74399286106 
    (index==692) ? 32'h3f3ead6e : // 0.7448338375 
    (index==693) ? 32'h3f3ee483 : // 0.745674324002 
    (index==694) ? 32'h3f3f1b90 : // 0.746514321138 
    (index==695) ? 32'h3f3f5294 : // 0.747353829478 
    (index==696) ? 32'h3f3f8991 : // 0.748192849589 
    (index==697) ? 32'h3f3fc085 : // 0.74903138204 
    (index==698) ? 32'h3f3ff771 : // 0.749869427397 
    (index==699) ? 32'h3f402e55 : // 0.750706986225 
    (index==700) ? 32'h3f406531 : // 0.751544059089 
    (index==701) ? 32'h3f409c04 : // 0.752380646553 
    (index==702) ? 32'h3f40d2d0 : // 0.753216749179 
    (index==703) ? 32'h3f410993 : // 0.754052367529 
    (index==704) ? 32'h3f41404e : // 0.754887502163 
    (index==705) ? 32'h3f417701 : // 0.755722153642 
    (index==706) ? 32'h3f41adac : // 0.756556322524 
    (index==707) ? 32'h3f41e44f : // 0.757390009367 
    (index==708) ? 32'h3f421aea : // 0.758223214727 
    (index==709) ? 32'h3f42517d : // 0.75905593916 
    (index==710) ? 32'h3f428808 : // 0.759888183222 
    (index==711) ? 32'h3f42be8a : // 0.760719947466 
    (index==712) ? 32'h3f42f505 : // 0.761551232444 
    (index==713) ? 32'h3f432b78 : // 0.76238203871 
    (index==714) ? 32'h3f4361e2 : // 0.763212366814 
    (index==715) ? 32'h3f439845 : // 0.764042217307 
    (index==716) ? 32'h3f43ce9f : // 0.764871590736 
    (index==717) ? 32'h3f4404f2 : // 0.765700487651 
    (index==718) ? 32'h3f443b3d : // 0.766528908599 
    (index==719) ? 32'h3f44717f : // 0.767356854126 
    (index==720) ? 32'h3f44a7ba : // 0.768184324777 
    (index==721) ? 32'h3f44dded : // 0.769011321097 
    (index==722) ? 32'h3f451417 : // 0.769837843629 
    (index==723) ? 32'h3f454a3a : // 0.770663892917 
    (index==724) ? 32'h3f458055 : // 0.771489469501 
    (index==725) ? 32'h3f45b668 : // 0.772314573922 
    (index==726) ? 32'h3f45ec73 : // 0.77313920672 
    (index==727) ? 32'h3f462276 : // 0.773963368434 
    (index==728) ? 32'h3f465871 : // 0.774787059601 
    (index==729) ? 32'h3f468e65 : // 0.77561028076 
    (index==730) ? 32'h3f46c450 : // 0.776433032445 
    (index==731) ? 32'h3f46fa34 : // 0.777255315192 
    (index==732) ? 32'h3f473010 : // 0.778077129535 
    (index==733) ? 32'h3f4765e3 : // 0.778898476008 
    (index==734) ? 32'h3f479bb0 : // 0.779719355143 
    (index==735) ? 32'h3f47d174 : // 0.780539767472 
    (index==736) ? 32'h3f480730 : // 0.781359713525 
    (index==737) ? 32'h3f483ce5 : // 0.782179193831 
    (index==738) ? 32'h3f487292 : // 0.78299820892 
    (index==739) ? 32'h3f48a837 : // 0.78381675932 
    (index==740) ? 32'h3f48ddd4 : // 0.784634845558 
    (index==741) ? 32'h3f491369 : // 0.785452468159 
    (index==742) ? 32'h3f4948f7 : // 0.786269627648 
    (index==743) ? 32'h3f497e7d : // 0.787086324552 
    (index==744) ? 32'h3f49b3fb : // 0.787902559391 
    (index==745) ? 32'h3f49e971 : // 0.78871833269 
    (index==746) ? 32'h3f4a1ee0 : // 0.78953364497 
    (index==747) ? 32'h3f4a5447 : // 0.790348496752 
    (index==748) ? 32'h3f4a89a6 : // 0.791162888555 
    (index==749) ? 32'h3f4abefe : // 0.791976820899 
    (index==750) ? 32'h3f4af44e : // 0.792790294301 
    (index==751) ? 32'h3f4b2996 : // 0.793603309279 
    (index==752) ? 32'h3f4b5ed6 : // 0.79441586635 
    (index==753) ? 32'h3f4b940f : // 0.795227966029 
    (index==754) ? 32'h3f4bc940 : // 0.79603960883 
    (index==755) ? 32'h3f4bfe69 : // 0.796850795267 
    (index==756) ? 32'h3f4c338b : // 0.797661525854 
    (index==757) ? 32'h3f4c68a5 : // 0.798471801102 
    (index==758) ? 32'h3f4c9db8 : // 0.799281621522 
    (index==759) ? 32'h3f4cd2c3 : // 0.800090987625 
    (index==760) ? 32'h3f4d07c6 : // 0.80089989992 
    (index==761) ? 32'h3f4d3cc2 : // 0.801708358916 
    (index==762) ? 32'h3f4d71b6 : // 0.802516365121 
    (index==763) ? 32'h3f4da6a2 : // 0.803323919041 
    (index==764) ? 32'h3f4ddb87 : // 0.804131021183 
    (index==765) ? 32'h3f4e1065 : // 0.804937672052 
    (index==766) ? 32'h3f4e453a : // 0.805743872152 
    (index==767) ? 32'h3f4e7a09 : // 0.806549621986 
    (index==768) ? 32'h3f4eaecf : // 0.807354922058 
    (index==769) ? 32'h3f4ee38f : // 0.808159772868 
    (index==770) ? 32'h3f4f1846 : // 0.808964174919 
    (index==771) ? 32'h3f4f4cf6 : // 0.80976812871 
    (index==772) ? 32'h3f4f819f : // 0.810571634741 
    (index==773) ? 32'h3f4fb640 : // 0.81137469351 
    (index==774) ? 32'h3f4feada : // 0.812177305514 
    (index==775) ? 32'h3f501f6c : // 0.812979471251 
    (index==776) ? 32'h3f5053f6 : // 0.813781191217 
    (index==777) ? 32'h3f508879 : // 0.814582465906 
    (index==778) ? 32'h3f50bcf5 : // 0.815383295814 
    (index==779) ? 32'h3f50f169 : // 0.816183681432 
    (index==780) ? 32'h3f5125d6 : // 0.816983623255 
    (index==781) ? 32'h3f515a3c : // 0.817783121775 
    (index==782) ? 32'h3f518e9a : // 0.818582177481 
    (index==783) ? 32'h3f51c2f0 : // 0.819380790865 
    (index==784) ? 32'h3f51f73f : // 0.820178962415 
    (index==785) ? 32'h3f522b87 : // 0.820976692621 
    (index==786) ? 32'h3f525fc7 : // 0.821773981971 
    (index==787) ? 32'h3f529400 : // 0.82257083095 
    (index==788) ? 32'h3f52c832 : // 0.823367240046 
    (index==789) ? 32'h3f52fc5c : // 0.824163209744 
    (index==790) ? 32'h3f53307e : // 0.824958740529 
    (index==791) ? 32'h3f53649a : // 0.825753832883 
    (index==792) ? 32'h3f5398ae : // 0.826548487291 
    (index==793) ? 32'h3f53ccbb : // 0.827342704234 
    (index==794) ? 32'h3f5400c0 : // 0.828136484194 
    (index==795) ? 32'h3f5434be : // 0.828929827651 
    (index==796) ? 32'h3f5468b5 : // 0.829722735086 
    (index==797) ? 32'h3f549ca5 : // 0.830515206977 
    (index==798) ? 32'h3f54d08d : // 0.831307243802 
    (index==799) ? 32'h3f55046e : // 0.832098846039 
    (index==800) ? 32'h3f553847 : // 0.832890014165 
    (index==801) ? 32'h3f556c19 : // 0.833680748655 
    (index==802) ? 32'h3f559fe5 : // 0.834471049984 
    (index==803) ? 32'h3f55d3a8 : // 0.835260918627 
    (index==804) ? 32'h3f560765 : // 0.836050355058 
    (index==805) ? 32'h3f563b1a : // 0.836839359749 
    (index==806) ? 32'h3f566ec8 : // 0.837627933171 
    (index==807) ? 32'h3f56a26f : // 0.838416075797 
    (index==808) ? 32'h3f56d60f : // 0.839203788097 
    (index==809) ? 32'h3f5709a7 : // 0.83999107054 
    (index==810) ? 32'h3f573d38 : // 0.840777923595 
    (index==811) ? 32'h3f5770c2 : // 0.841564347731 
    (index==812) ? 32'h3f57a445 : // 0.842350343414 
    (index==813) ? 32'h3f57d7c1 : // 0.843135911111 
    (index==814) ? 32'h3f580b35 : // 0.843921051289 
    (index==815) ? 32'h3f583ea3 : // 0.844705764412 
    (index==816) ? 32'h3f587209 : // 0.845490050944 
    (index==817) ? 32'h3f58a568 : // 0.84627391135 
    (index==818) ? 32'h3f58d8c0 : // 0.847057346091 
    (index==819) ? 32'h3f590c10 : // 0.847840355631 
    (index==820) ? 32'h3f593f5a : // 0.848622940429 
    (index==821) ? 32'h3f59729c : // 0.849405100948 
    (index==822) ? 32'h3f59a5d8 : // 0.850186837646 
    (index==823) ? 32'h3f59d90c : // 0.850968150982 
    (index==824) ? 32'h3f5a0c39 : // 0.851749041416 
    (index==825) ? 32'h3f5a3f5f : // 0.852529509404 
    (index==826) ? 32'h3f5a727e : // 0.853309555404 
    (index==827) ? 32'h3f5aa596 : // 0.854089179871 
    (index==828) ? 32'h3f5ad8a7 : // 0.85486838326 
    (index==829) ? 32'h3f5b0bb1 : // 0.855647166027 
    (index==830) ? 32'h3f5b3eb4 : // 0.856425528626 
    (index==831) ? 32'h3f5b71af : // 0.857203471508 
    (index==832) ? 32'h3f5ba4a4 : // 0.857980995128 
    (index==833) ? 32'h3f5bd792 : // 0.858758099935 
    (index==834) ? 32'h3f5c0a78 : // 0.859534786383 
    (index==835) ? 32'h3f5c3d58 : // 0.860311054919 
    (index==836) ? 32'h3f5c7031 : // 0.861086905995 
    (index==837) ? 32'h3f5ca302 : // 0.861862340059 
    (index==838) ? 32'h3f5cd5cd : // 0.862637357559 
    (index==839) ? 32'h3f5d0890 : // 0.863411958942 
    (index==840) ? 32'h3f5d3b4d : // 0.864186144654 
    (index==841) ? 32'h3f5d6e03 : // 0.864959915143 
    (index==842) ? 32'h3f5da0b2 : // 0.865733270852 
    (index==843) ? 32'h3f5dd359 : // 0.866506212226 
    (index==844) ? 32'h3f5e05fa : // 0.86727873971 
    (index==845) ? 32'h3f5e3894 : // 0.868050853745 
    (index==846) ? 32'h3f5e6b27 : // 0.868822554775 
    (index==847) ? 32'h3f5e9db3 : // 0.869593843241 
    (index==848) ? 32'h3f5ed038 : // 0.870364719583 
    (index==849) ? 32'h3f5f02b7 : // 0.871135184243 
    (index==850) ? 32'h3f5f352e : // 0.871905237659 
    (index==851) ? 32'h3f5f679e : // 0.872674880271 
    (index==852) ? 32'h3f5f9a08 : // 0.873444112515 
    (index==853) ? 32'h3f5fcc6b : // 0.874212934831 
    (index==854) ? 32'h3f5ffec7 : // 0.874981347654 
    (index==855) ? 32'h3f60311c : // 0.87574935142 
    (index==856) ? 32'h3f60636a : // 0.876516946565 
    (index==857) ? 32'h3f6095b1 : // 0.877284133523 
    (index==858) ? 32'h3f60c7f1 : // 0.878050912729 
    (index==859) ? 32'h3f60fa2b : // 0.878817284614 
    (index==860) ? 32'h3f612c5e : // 0.879583249613 
    (index==861) ? 32'h3f615e8a : // 0.880348808156 
    (index==862) ? 32'h3f6190af : // 0.881113960675 
    (index==863) ? 32'h3f61c2cd : // 0.8818787076 
    (index==864) ? 32'h3f61f4e5 : // 0.882643049362 
    (index==865) ? 32'h3f6226f5 : // 0.883406986388 
    (index==866) ? 32'h3f6258ff : // 0.884170519108 
    (index==867) ? 32'h3f628b02 : // 0.88493364795 
    (index==868) ? 32'h3f62bcff : // 0.885696373339 
    (index==869) ? 32'h3f62eef5 : // 0.886458695704 
    (index==870) ? 32'h3f6320e3 : // 0.887220615468 
    (index==871) ? 32'h3f6352cc : // 0.887982133058 
    (index==872) ? 32'h3f6384ad : // 0.888743248898 
    (index==873) ? 32'h3f63b688 : // 0.889503963411 
    (index==874) ? 32'h3f63e85c : // 0.890264277021 
    (index==875) ? 32'h3f641a29 : // 0.891024190149 
    (index==876) ? 32'h3f644bef : // 0.891783703218 
    (index==877) ? 32'h3f647daf : // 0.892542816649 
    (index==878) ? 32'h3f64af68 : // 0.893301530861 
    (index==879) ? 32'h3f64e11b : // 0.894059846274 
    (index==880) ? 32'h3f6512c6 : // 0.894817763308 
    (index==881) ? 32'h3f65446b : // 0.895575282381 
    (index==882) ? 32'h3f65760a : // 0.89633240391 
    (index==883) ? 32'h3f65a7a2 : // 0.897089128313 
    (index==884) ? 32'h3f65d933 : // 0.897845456006 
    (index==885) ? 32'h3f660abd : // 0.898601387404 
    (index==886) ? 32'h3f663c41 : // 0.899356922923 
    (index==887) ? 32'h3f666dbe : // 0.900112062977 
    (index==888) ? 32'h3f669f35 : // 0.900866807981 
    (index==889) ? 32'h3f66d0a4 : // 0.901621158346 
    (index==890) ? 32'h3f67020e : // 0.902375114486 
    (index==891) ? 32'h3f673370 : // 0.903128676812 
    (index==892) ? 32'h3f6764cc : // 0.903881845736 
    (index==893) ? 32'h3f679622 : // 0.904634621668 
    (index==894) ? 32'h3f67c771 : // 0.905387005018 
    (index==895) ? 32'h3f67f8b9 : // 0.906138996195 
    (index==896) ? 32'h3f6829fb : // 0.906890595609 
    (index==897) ? 32'h3f685b36 : // 0.907641803666 
    (index==898) ? 32'h3f688c6b : // 0.908392620774 
    (index==899) ? 32'h3f68bd99 : // 0.90914304734 
    (index==900) ? 32'h3f68eec0 : // 0.90989308377 
    (index==901) ? 32'h3f691fe1 : // 0.91064273047 
    (index==902) ? 32'h3f6950fc : // 0.911391987843 
    (index==903) ? 32'h3f698210 : // 0.912140856296 
    (index==904) ? 32'h3f69b31d : // 0.91288933623 
    (index==905) ? 32'h3f69e424 : // 0.913637428049 
    (index==906) ? 32'h3f6a1524 : // 0.914385132155 
    (index==907) ? 32'h3f6a461e : // 0.915132448951 
    (index==908) ? 32'h3f6a7712 : // 0.915879378836 
    (index==909) ? 32'h3f6aa7ff : // 0.916625922211 
    (index==910) ? 32'h3f6ad8e5 : // 0.917372079477 
    (index==911) ? 32'h3f6b09c5 : // 0.918117851032 
    (index==912) ? 32'h3f6b3a9f : // 0.918863237275 
    (index==913) ? 32'h3f6b6b72 : // 0.919608238603 
    (index==914) ? 32'h3f6b9c3e : // 0.920352855415 
    (index==915) ? 32'h3f6bcd04 : // 0.921097088107 
    (index==916) ? 32'h3f6bfdc4 : // 0.921840937074 
    (index==917) ? 32'h3f6c2e7d : // 0.922584402714 
    (index==918) ? 32'h3f6c5f30 : // 0.923327485419 
    (index==919) ? 32'h3f6c8fdd : // 0.924070185585 
    (index==920) ? 32'h3f6cc083 : // 0.924812503606 
    (index==921) ? 32'h3f6cf122 : // 0.925554439874 
    (index==922) ? 32'h3f6d21bb : // 0.926295994781 
    (index==923) ? 32'h3f6d524e : // 0.92703716872 
    (index==924) ? 32'h3f6d82db : // 0.927777962082 
    (index==925) ? 32'h3f6db361 : // 0.928518375258 
    (index==926) ? 32'h3f6de3e1 : // 0.929258408637 
    (index==927) ? 32'h3f6e145a : // 0.929998062609 
    (index==928) ? 32'h3f6e44cd : // 0.930737337563 
    (index==929) ? 32'h3f6e7539 : // 0.931476233887 
    (index==930) ? 32'h3f6ea5a0 : // 0.932214751968 
    (index==931) ? 32'h3f6ed600 : // 0.932952892195 
    (index==932) ? 32'h3f6f0659 : // 0.933690654952 
    (index==933) ? 32'h3f6f36ad : // 0.934428040627 
    (index==934) ? 32'h3f6f66fa : // 0.935165049604 
    (index==935) ? 32'h3f6f9740 : // 0.935901682268 
    (index==936) ? 32'h3f6fc781 : // 0.936637939003 
    (index==937) ? 32'h3f6ff7bb : // 0.937373820192 
    (index==938) ? 32'h3f7027ee : // 0.938109326219 
    (index==939) ? 32'h3f70581c : // 0.938844457466 
    (index==940) ? 32'h3f708843 : // 0.939579214315 
    (index==941) ? 32'h3f70b864 : // 0.940313597146 
    (index==942) ? 32'h3f70e87e : // 0.941047606341 
    (index==943) ? 32'h3f711893 : // 0.941781242279 
    (index==944) ? 32'h3f7148a1 : // 0.942514505339 
    (index==945) ? 32'h3f7178a9 : // 0.943247395902 
    (index==946) ? 32'h3f71a8aa : // 0.943979914344 
    (index==947) ? 32'h3f71d8a6 : // 0.944712061043 
    (index==948) ? 32'h3f72089b : // 0.945443836378 
    (index==949) ? 32'h3f72388a : // 0.946175240724 
    (index==950) ? 32'h3f726873 : // 0.946906274456 
    (index==951) ? 32'h3f729855 : // 0.947636937952 
    (index==952) ? 32'h3f72c831 : // 0.948367231585 
    (index==953) ? 32'h3f72f807 : // 0.949097155729 
    (index==954) ? 32'h3f7327d7 : // 0.949826710759 
    (index==955) ? 32'h3f7357a1 : // 0.950555897048 
    (index==956) ? 32'h3f738765 : // 0.951284714967 
    (index==957) ? 32'h3f73b722 : // 0.952013164889 
    (index==958) ? 32'h3f73e6d9 : // 0.952741247186 
    (index==959) ? 32'h3f74168a : // 0.953468962229 
    (index==960) ? 32'h3f744635 : // 0.954196310387 
    (index==961) ? 32'h3f7475da : // 0.95492329203 
    (index==962) ? 32'h3f74a578 : // 0.955649907528 
    (index==963) ? 32'h3f74d511 : // 0.95637615725 
    (index==964) ? 32'h3f7504a3 : // 0.957102041562 
    (index==965) ? 32'h3f75342f : // 0.957827560834 
    (index==966) ? 32'h3f7563b5 : // 0.958552715431 
    (index==967) ? 32'h3f759335 : // 0.959277505721 
    (index==968) ? 32'h3f75c2af : // 0.960001932068 
    (index==969) ? 32'h3f75f223 : // 0.960725994839 
    (index==970) ? 32'h3f762191 : // 0.961449694398 
    (index==971) ? 32'h3f7650f8 : // 0.96217303111 
    (index==972) ? 32'h3f76805a : // 0.962896005337 
    (index==973) ? 32'h3f76afb5 : // 0.963618617444 
    (index==974) ? 32'h3f76df0b : // 0.964340867792 
    (index==975) ? 32'h3f770e5a : // 0.965062756745 
    (index==976) ? 32'h3f773da3 : // 0.965784284662 
    (index==977) ? 32'h3f776ce6 : // 0.966505451906 
    (index==978) ? 32'h3f779c23 : // 0.967226258836 
    (index==979) ? 32'h3f77cb5a : // 0.967946705813 
    (index==980) ? 32'h3f77fa8c : // 0.968666793195 
    (index==981) ? 32'h3f7829b7 : // 0.969386521342 
    (index==982) ? 32'h3f7858dc : // 0.970105890612 
    (index==983) ? 32'h3f7887fb : // 0.970824901363 
    (index==984) ? 32'h3f78b714 : // 0.971543553951 
    (index==985) ? 32'h3f78e627 : // 0.972261848733 
    (index==986) ? 32'h3f791534 : // 0.972979786066 
    (index==987) ? 32'h3f79443b : // 0.973697366305 
    (index==988) ? 32'h3f79733c : // 0.974414589806 
    (index==989) ? 32'h3f79a237 : // 0.975131456921 
    (index==990) ? 32'h3f79d12c : // 0.975847968007 
    (index==991) ? 32'h3f7a001b : // 0.976564123415 
    (index==992) ? 32'h3f7a2f04 : // 0.9772799235 
    (index==993) ? 32'h3f7a5de7 : // 0.977995368613 
    (index==994) ? 32'h3f7a8cc4 : // 0.978710459106 
    (index==995) ? 32'h3f7abb9c : // 0.979425195331 
    (index==996) ? 32'h3f7aea6d : // 0.980139577639 
    (index==997) ? 32'h3f7b1938 : // 0.98085360638 
    (index==998) ? 32'h3f7b47fe : // 0.981567281903 
    (index==999) ? 32'h3f7b76bd : // 0.982280604558 
    (index==1000) ? 32'h3f7ba577 : // 0.982993574694 
    (index==1001) ? 32'h3f7bd42b : // 0.983706192659 
    (index==1002) ? 32'h3f7c02d9 : // 0.984418458801 
    (index==1003) ? 32'h3f7c3181 : // 0.985130373467 
    (index==1004) ? 32'h3f7c6023 : // 0.985841937003 
    (index==1005) ? 32'h3f7c8ebf : // 0.986553149757 
    (index==1006) ? 32'h3f7cbd55 : // 0.987264012073 
    (index==1007) ? 32'h3f7cebe5 : // 0.987974524296 
    (index==1008) ? 32'h3f7d1a70 : // 0.988684686772 
    (index==1009) ? 32'h3f7d48f5 : // 0.989394499845 
    (index==1010) ? 32'h3f7d7774 : // 0.990103963858 
    (index==1011) ? 32'h3f7da5ed : // 0.990813079154 
    (index==1012) ? 32'h3f7dd460 : // 0.991521846076 
    (index==1013) ? 32'h3f7e02cd : // 0.992230264966 
    (index==1014) ? 32'h3f7e3134 : // 0.992938336166 
    (index==1015) ? 32'h3f7e5f96 : // 0.993646060017 
    (index==1016) ? 32'h3f7e8df2 : // 0.994353436859 
    (index==1017) ? 32'h3f7ebc48 : // 0.995060467033 
    (index==1018) ? 32'h3f7eea98 : // 0.995767150878 
    (index==1019) ? 32'h3f7f18e2 : // 0.996473488733 
    (index==1020) ? 32'h3f7f4727 : // 0.997179480938 
    (index==1021) ? 32'h3f7f7566 : // 0.997885127829 
    (index==1022) ? 32'h3f7fa39f : // 0.998590429745 
    (index==1023) ? 32'h3f7fd1d2 : // 0.999295387023 
    0;
endmodule
