module atan_table_till_2(input [9:0] addr,output [24:0] result,output [24:0] lastone);
 // tablesize = 1024
assign result = 
    (addr==0) ? 0 :  //   in=0.000000 val=0.000000
    (addr==1) ? 32767 :  //   in=0.001953 val=0.001953
    (addr==2) ? 65535 :  //   in=0.003906 val=0.003906
    (addr==3) ? 98302 :  //   in=0.005859 val=0.005859
    (addr==4) ? 131069 :  //   in=0.007812 val=0.007812
    (addr==5) ? 163834 :  //   in=0.009766 val=0.009765
    (addr==6) ? 196599 :  //   in=0.011719 val=0.011718
    (addr==7) ? 229361 :  //   in=0.013672 val=0.013671
    (addr==8) ? 262122 :  //   in=0.015625 val=0.015624
    (addr==9) ? 294881 :  //   in=0.017578 val=0.017576
    (addr==10) ? 327638 :  //   in=0.019531 val=0.019529
    (addr==11) ? 360392 :  //   in=0.021484 val=0.021481
    (addr==12) ? 393144 :  //   in=0.023438 val=0.023433
    (addr==13) ? 425892 :  //   in=0.025391 val=0.025385
    (addr==14) ? 458637 :  //   in=0.027344 val=0.027337
    (addr==15) ? 491379 :  //   in=0.029297 val=0.029288
    (addr==16) ? 524117 :  //   in=0.031250 val=0.031240
    (addr==17) ? 556851 :  //   in=0.033203 val=0.033191
    (addr==18) ? 589581 :  //   in=0.035156 val=0.035142
    (addr==19) ? 622306 :  //   in=0.037109 val=0.037092
    (addr==20) ? 655026 :  //   in=0.039062 val=0.039043
    (addr==21) ? 687742 :  //   in=0.041016 val=0.040993
    (addr==22) ? 720452 :  //   in=0.042969 val=0.042942
    (addr==23) ? 753157 :  //   in=0.044922 val=0.044892
    (addr==24) ? 785856 :  //   in=0.046875 val=0.046841
    (addr==25) ? 818549 :  //   in=0.048828 val=0.048789
    (addr==26) ? 851236 :  //   in=0.050781 val=0.050738
    (addr==27) ? 883917 :  //   in=0.052734 val=0.052686
    (addr==28) ? 916590 :  //   in=0.054688 val=0.054633
    (addr==29) ? 949257 :  //   in=0.056641 val=0.056580
    (addr==30) ? 981917 :  //   in=0.058594 val=0.058527
    (addr==31) ? 1014569 :  //   in=0.060547 val=0.060473
    (addr==32) ? 1047213 :  //   in=0.062500 val=0.062419
    (addr==33) ? 1079850 :  //   in=0.064453 val=0.064364
    (addr==34) ? 1112478 :  //   in=0.066406 val=0.066309
    (addr==35) ? 1145098 :  //   in=0.068359 val=0.068253
    (addr==36) ? 1177709 :  //   in=0.070312 val=0.070197
    (addr==37) ? 1210312 :  //   in=0.072266 val=0.072140
    (addr==38) ? 1242905 :  //   in=0.074219 val=0.074083
    (addr==39) ? 1275488 :  //   in=0.076172 val=0.076025
    (addr==40) ? 1308063 :  //   in=0.078125 val=0.077967
    (addr==41) ? 1340627 :  //   in=0.080078 val=0.079908
    (addr==42) ? 1373181 :  //   in=0.082031 val=0.081848
    (addr==43) ? 1405725 :  //   in=0.083984 val=0.083788
    (addr==44) ? 1438258 :  //   in=0.085938 val=0.085727
    (addr==45) ? 1470780 :  //   in=0.087891 val=0.087665
    (addr==46) ? 1503291 :  //   in=0.089844 val=0.089603
    (addr==47) ? 1535791 :  //   in=0.091797 val=0.091540
    (addr==48) ? 1568280 :  //   in=0.093750 val=0.093477
    (addr==49) ? 1600756 :  //   in=0.095703 val=0.095413
    (addr==50) ? 1633221 :  //   in=0.097656 val=0.097348
    (addr==51) ? 1665673 :  //   in=0.099609 val=0.099282
    (addr==52) ? 1698113 :  //   in=0.101562 val=0.101215
    (addr==53) ? 1730540 :  //   in=0.103516 val=0.103148
    (addr==54) ? 1762954 :  //   in=0.105469 val=0.105080
    (addr==55) ? 1795355 :  //   in=0.107422 val=0.107012
    (addr==56) ? 1827742 :  //   in=0.109375 val=0.108942
    (addr==57) ? 1860116 :  //   in=0.111328 val=0.110872
    (addr==58) ? 1892476 :  //   in=0.113281 val=0.112800
    (addr==59) ? 1924822 :  //   in=0.115234 val=0.114728
    (addr==60) ? 1957153 :  //   in=0.117188 val=0.116655
    (addr==61) ? 1989470 :  //   in=0.119141 val=0.118582
    (addr==62) ? 2021772 :  //   in=0.121094 val=0.120507
    (addr==63) ? 2054059 :  //   in=0.123047 val=0.122431
    (addr==64) ? 2086330 :  //   in=0.125000 val=0.124355
    (addr==65) ? 2118586 :  //   in=0.126953 val=0.126278
    (addr==66) ? 2150827 :  //   in=0.128906 val=0.128199
    (addr==67) ? 2183051 :  //   in=0.130859 val=0.130120
    (addr==68) ? 2215259 :  //   in=0.132812 val=0.132040
    (addr==69) ? 2247451 :  //   in=0.134766 val=0.133959
    (addr==70) ? 2279626 :  //   in=0.136719 val=0.135876
    (addr==71) ? 2311784 :  //   in=0.138672 val=0.137793
    (addr==72) ? 2343925 :  //   in=0.140625 val=0.139709
    (addr==73) ? 2376049 :  //   in=0.142578 val=0.141624
    (addr==74) ? 2408156 :  //   in=0.144531 val=0.143537
    (addr==75) ? 2440244 :  //   in=0.146484 val=0.145450
    (addr==76) ? 2472315 :  //   in=0.148438 val=0.147361
    (addr==77) ? 2504367 :  //   in=0.150391 val=0.149272
    (addr==78) ? 2536401 :  //   in=0.152344 val=0.151181
    (addr==79) ? 2568417 :  //   in=0.154297 val=0.153090
    (addr==80) ? 2600413 :  //   in=0.156250 val=0.154997
    (addr==81) ? 2632391 :  //   in=0.158203 val=0.156903
    (addr==82) ? 2664349 :  //   in=0.160156 val=0.158808
    (addr==83) ? 2696288 :  //   in=0.162109 val=0.160711
    (addr==84) ? 2728207 :  //   in=0.164062 val=0.162614
    (addr==85) ? 2760106 :  //   in=0.166016 val=0.164515
    (addr==86) ? 2791985 :  //   in=0.167969 val=0.166415
    (addr==87) ? 2823844 :  //   in=0.169922 val=0.168314
    (addr==88) ? 2855682 :  //   in=0.171875 val=0.170212
    (addr==89) ? 2887499 :  //   in=0.173828 val=0.172108
    (addr==90) ? 2919295 :  //   in=0.175781 val=0.174004
    (addr==91) ? 2951071 :  //   in=0.177734 val=0.175898
    (addr==92) ? 2982825 :  //   in=0.179688 val=0.177790
    (addr==93) ? 3014557 :  //   in=0.181641 val=0.179682
    (addr==94) ? 3046267 :  //   in=0.183594 val=0.181572
    (addr==95) ? 3077956 :  //   in=0.185547 val=0.183460
    (addr==96) ? 3109622 :  //   in=0.187500 val=0.185348
    (addr==97) ? 3141266 :  //   in=0.189453 val=0.187234
    (addr==98) ? 3172887 :  //   in=0.191406 val=0.189119
    (addr==99) ? 3204486 :  //   in=0.193359 val=0.191002
    (addr==100) ? 3236061 :  //   in=0.195312 val=0.192884
    (addr==101) ? 3267614 :  //   in=0.197266 val=0.194765
    (addr==102) ? 3299142 :  //   in=0.199219 val=0.196644
    (addr==103) ? 3330648 :  //   in=0.201172 val=0.198522
    (addr==104) ? 3362129 :  //   in=0.203125 val=0.200399
    (addr==105) ? 3393587 :  //   in=0.205078 val=0.202274
    (addr==106) ? 3425020 :  //   in=0.207031 val=0.204147
    (addr==107) ? 3456429 :  //   in=0.208984 val=0.206019
    (addr==108) ? 3487814 :  //   in=0.210938 val=0.207890
    (addr==109) ? 3519173 :  //   in=0.212891 val=0.209759
    (addr==110) ? 3550508 :  //   in=0.214844 val=0.211627
    (addr==111) ? 3581818 :  //   in=0.216797 val=0.213493
    (addr==112) ? 3613102 :  //   in=0.218750 val=0.215358
    (addr==113) ? 3644361 :  //   in=0.220703 val=0.217221
    (addr==114) ? 3675594 :  //   in=0.222656 val=0.219083
    (addr==115) ? 3706801 :  //   in=0.224609 val=0.220943
    (addr==116) ? 3737983 :  //   in=0.226562 val=0.222801
    (addr==117) ? 3769138 :  //   in=0.228516 val=0.224658
    (addr==118) ? 3800266 :  //   in=0.230469 val=0.226514
    (addr==119) ? 3831368 :  //   in=0.232422 val=0.228367
    (addr==120) ? 3862443 :  //   in=0.234375 val=0.230220
    (addr==121) ? 3893491 :  //   in=0.236328 val=0.232070
    (addr==122) ? 3924513 :  //   in=0.238281 val=0.233919
    (addr==123) ? 3955506 :  //   in=0.240234 val=0.235767
    (addr==124) ? 3986473 :  //   in=0.242188 val=0.237612
    (addr==125) ? 4017411 :  //   in=0.244141 val=0.239456
    (addr==126) ? 4048322 :  //   in=0.246094 val=0.241299
    (addr==127) ? 4079205 :  //   in=0.248047 val=0.243140
    (addr==128) ? 4110059 :  //   in=0.250000 val=0.244979
    (addr==129) ? 4140886 :  //   in=0.251953 val=0.246816
    (addr==130) ? 4171683 :  //   in=0.253906 val=0.248652
    (addr==131) ? 4202453 :  //   in=0.255859 val=0.250486
    (addr==132) ? 4233193 :  //   in=0.257812 val=0.252318
    (addr==133) ? 4263904 :  //   in=0.259766 val=0.254149
    (addr==134) ? 4294586 :  //   in=0.261719 val=0.255977
    (addr==135) ? 4325239 :  //   in=0.263672 val=0.257804
    (addr==136) ? 4355862 :  //   in=0.265625 val=0.259630
    (addr==137) ? 4386455 :  //   in=0.267578 val=0.261453
    (addr==138) ? 4417019 :  //   in=0.269531 val=0.263275
    (addr==139) ? 4447553 :  //   in=0.271484 val=0.265095
    (addr==140) ? 4478056 :  //   in=0.273438 val=0.266913
    (addr==141) ? 4508530 :  //   in=0.275391 val=0.268729
    (addr==142) ? 4538972 :  //   in=0.277344 val=0.270544
    (addr==143) ? 4569385 :  //   in=0.279297 val=0.272357
    (addr==144) ? 4599766 :  //   in=0.281250 val=0.274167
    (addr==145) ? 4630117 :  //   in=0.283203 val=0.275976
    (addr==146) ? 4660436 :  //   in=0.285156 val=0.277784
    (addr==147) ? 4690724 :  //   in=0.287109 val=0.279589
    (addr==148) ? 4720981 :  //   in=0.289062 val=0.281392
    (addr==149) ? 4751206 :  //   in=0.291016 val=0.283194
    (addr==150) ? 4781400 :  //   in=0.292969 val=0.284994
    (addr==151) ? 4811562 :  //   in=0.294922 val=0.286791
    (addr==152) ? 4841692 :  //   in=0.296875 val=0.288587
    (addr==153) ? 4871790 :  //   in=0.298828 val=0.290381
    (addr==154) ? 4901855 :  //   in=0.300781 val=0.292173
    (addr==155) ? 4931889 :  //   in=0.302734 val=0.293964
    (addr==156) ? 4961889 :  //   in=0.304688 val=0.295752
    (addr==157) ? 4991857 :  //   in=0.306641 val=0.297538
    (addr==158) ? 5021793 :  //   in=0.308594 val=0.299322
    (addr==159) ? 5051695 :  //   in=0.310547 val=0.301105
    (addr==160) ? 5081564 :  //   in=0.312500 val=0.302885
    (addr==161) ? 5111400 :  //   in=0.314453 val=0.304663
    (addr==162) ? 5141203 :  //   in=0.316406 val=0.306440
    (addr==163) ? 5170972 :  //   in=0.318359 val=0.308214
    (addr==164) ? 5200708 :  //   in=0.320312 val=0.309986
    (addr==165) ? 5230410 :  //   in=0.322266 val=0.311757
    (addr==166) ? 5260078 :  //   in=0.324219 val=0.313525
    (addr==167) ? 5289712 :  //   in=0.326172 val=0.315291
    (addr==168) ? 5319312 :  //   in=0.328125 val=0.317056
    (addr==169) ? 5348878 :  //   in=0.330078 val=0.318818
    (addr==170) ? 5378410 :  //   in=0.332031 val=0.320578
    (addr==171) ? 5407907 :  //   in=0.333984 val=0.322336
    (addr==172) ? 5437369 :  //   in=0.335938 val=0.324092
    (addr==173) ? 5466797 :  //   in=0.337891 val=0.325846
    (addr==174) ? 5496189 :  //   in=0.339844 val=0.327598
    (addr==175) ? 5525547 :  //   in=0.341797 val=0.329348
    (addr==176) ? 5554870 :  //   in=0.343750 val=0.331096
    (addr==177) ? 5584157 :  //   in=0.345703 val=0.332842
    (addr==178) ? 5613410 :  //   in=0.347656 val=0.334585
    (addr==179) ? 5642627 :  //   in=0.349609 val=0.336327
    (addr==180) ? 5671808 :  //   in=0.351562 val=0.338066
    (addr==181) ? 5700954 :  //   in=0.353516 val=0.339803
    (addr==182) ? 5730063 :  //   in=0.355469 val=0.341538
    (addr==183) ? 5759137 :  //   in=0.357422 val=0.343271
    (addr==184) ? 5788176 :  //   in=0.359375 val=0.345002
    (addr==185) ? 5817178 :  //   in=0.361328 val=0.346731
    (addr==186) ? 5846143 :  //   in=0.363281 val=0.348457
    (addr==187) ? 5875073 :  //   in=0.365234 val=0.350182
    (addr==188) ? 5903966 :  //   in=0.367188 val=0.351904
    (addr==189) ? 5932823 :  //   in=0.369141 val=0.353624
    (addr==190) ? 5961643 :  //   in=0.371094 val=0.355342
    (addr==191) ? 5990426 :  //   in=0.373047 val=0.357057
    (addr==192) ? 6019173 :  //   in=0.375000 val=0.358771
    (addr==193) ? 6047882 :  //   in=0.376953 val=0.360482
    (addr==194) ? 6076555 :  //   in=0.378906 val=0.362191
    (addr==195) ? 6105190 :  //   in=0.380859 val=0.363898
    (addr==196) ? 6133789 :  //   in=0.382812 val=0.365602
    (addr==197) ? 6162350 :  //   in=0.384766 val=0.367305
    (addr==198) ? 6190874 :  //   in=0.386719 val=0.369005
    (addr==199) ? 6219360 :  //   in=0.388672 val=0.370703
    (addr==200) ? 6247809 :  //   in=0.390625 val=0.372398
    (addr==201) ? 6276220 :  //   in=0.392578 val=0.374092
    (addr==202) ? 6304593 :  //   in=0.394531 val=0.375783
    (addr==203) ? 6332929 :  //   in=0.396484 val=0.377472
    (addr==204) ? 6361226 :  //   in=0.398438 val=0.379159
    (addr==205) ? 6389486 :  //   in=0.400391 val=0.380843
    (addr==206) ? 6417708 :  //   in=0.402344 val=0.382525
    (addr==207) ? 6445891 :  //   in=0.404297 val=0.384205
    (addr==208) ? 6474036 :  //   in=0.406250 val=0.385883
    (addr==209) ? 6502143 :  //   in=0.408203 val=0.387558
    (addr==210) ? 6530212 :  //   in=0.410156 val=0.389231
    (addr==211) ? 6558242 :  //   in=0.412109 val=0.390902
    (addr==212) ? 6586233 :  //   in=0.414062 val=0.392570
    (addr==213) ? 6614186 :  //   in=0.416016 val=0.394236
    (addr==214) ? 6642101 :  //   in=0.417969 val=0.395900
    (addr==215) ? 6669976 :  //   in=0.419922 val=0.397562
    (addr==216) ? 6697813 :  //   in=0.421875 val=0.399221
    (addr==217) ? 6725610 :  //   in=0.423828 val=0.400878
    (addr==218) ? 6753369 :  //   in=0.425781 val=0.402532
    (addr==219) ? 6781089 :  //   in=0.427734 val=0.404184
    (addr==220) ? 6808769 :  //   in=0.429688 val=0.405834
    (addr==221) ? 6836410 :  //   in=0.431641 val=0.407482
    (addr==222) ? 6864012 :  //   in=0.433594 val=0.409127
    (addr==223) ? 6891575 :  //   in=0.435547 val=0.410770
    (addr==224) ? 6919099 :  //   in=0.437500 val=0.412410
    (addr==225) ? 6946582 :  //   in=0.439453 val=0.414049
    (addr==226) ? 6974027 :  //   in=0.441406 val=0.415684
    (addr==227) ? 7001432 :  //   in=0.443359 val=0.417318
    (addr==228) ? 7028797 :  //   in=0.445312 val=0.418949
    (addr==229) ? 7056122 :  //   in=0.447266 val=0.420578
    (addr==230) ? 7083408 :  //   in=0.449219 val=0.422204
    (addr==231) ? 7110654 :  //   in=0.451172 val=0.423828
    (addr==232) ? 7137860 :  //   in=0.453125 val=0.425450
    (addr==233) ? 7165026 :  //   in=0.455078 val=0.427069
    (addr==234) ? 7192152 :  //   in=0.457031 val=0.428686
    (addr==235) ? 7219238 :  //   in=0.458984 val=0.430300
    (addr==236) ? 7246284 :  //   in=0.460938 val=0.431912
    (addr==237) ? 7273290 :  //   in=0.462891 val=0.433522
    (addr==238) ? 7300256 :  //   in=0.464844 val=0.435129
    (addr==239) ? 7327181 :  //   in=0.466797 val=0.436734
    (addr==240) ? 7354067 :  //   in=0.468750 val=0.438337
    (addr==241) ? 7380912 :  //   in=0.470703 val=0.439937
    (addr==242) ? 7407716 :  //   in=0.472656 val=0.441534
    (addr==243) ? 7434480 :  //   in=0.474609 val=0.443130
    (addr==244) ? 7461204 :  //   in=0.476562 val=0.444722
    (addr==245) ? 7487887 :  //   in=0.478516 val=0.446313
    (addr==246) ? 7514529 :  //   in=0.480469 val=0.447901
    (addr==247) ? 7541131 :  //   in=0.482422 val=0.449486
    (addr==248) ? 7567693 :  //   in=0.484375 val=0.451070
    (addr==249) ? 7594213 :  //   in=0.486328 val=0.452650
    (addr==250) ? 7620693 :  //   in=0.488281 val=0.454229
    (addr==251) ? 7647132 :  //   in=0.490234 val=0.455805
    (addr==252) ? 7673531 :  //   in=0.492188 val=0.457378
    (addr==253) ? 7699888 :  //   in=0.494141 val=0.458949
    (addr==254) ? 7726205 :  //   in=0.496094 val=0.460518
    (addr==255) ? 7752481 :  //   in=0.498047 val=0.462084
    (addr==256) ? 7778716 :  //   in=0.500000 val=0.463648
    (addr==257) ? 7804909 :  //   in=0.501953 val=0.465209
    (addr==258) ? 7831062 :  //   in=0.503906 val=0.466768
    (addr==259) ? 7857174 :  //   in=0.505859 val=0.468324
    (addr==260) ? 7883245 :  //   in=0.507812 val=0.469878
    (addr==261) ? 7909275 :  //   in=0.509766 val=0.471430
    (addr==262) ? 7935264 :  //   in=0.511719 val=0.472979
    (addr==263) ? 7961211 :  //   in=0.513672 val=0.474525
    (addr==264) ? 7987117 :  //   in=0.515625 val=0.476069
    (addr==265) ? 8012983 :  //   in=0.517578 val=0.477611
    (addr==266) ? 8038807 :  //   in=0.519531 val=0.479150
    (addr==267) ? 8064589 :  //   in=0.521484 val=0.480687
    (addr==268) ? 8090331 :  //   in=0.523438 val=0.482221
    (addr==269) ? 8116031 :  //   in=0.525391 val=0.483753
    (addr==270) ? 8141690 :  //   in=0.527344 val=0.485283
    (addr==271) ? 8167307 :  //   in=0.529297 val=0.486809
    (addr==272) ? 8192884 :  //   in=0.531250 val=0.488334
    (addr==273) ? 8218419 :  //   in=0.533203 val=0.489856
    (addr==274) ? 8243912 :  //   in=0.535156 val=0.491375
    (addr==275) ? 8269364 :  //   in=0.537109 val=0.492893
    (addr==276) ? 8294775 :  //   in=0.539062 val=0.494407
    (addr==277) ? 8320144 :  //   in=0.541016 val=0.495919
    (addr==278) ? 8345472 :  //   in=0.542969 val=0.497429
    (addr==279) ? 8370758 :  //   in=0.544922 val=0.498936
    (addr==280) ? 8396003 :  //   in=0.546875 val=0.500441
    (addr==281) ? 8421207 :  //   in=0.548828 val=0.501943
    (addr==282) ? 8446368 :  //   in=0.550781 val=0.503443
    (addr==283) ? 8471489 :  //   in=0.552734 val=0.504940
    (addr==284) ? 8496568 :  //   in=0.554688 val=0.506435
    (addr==285) ? 8521605 :  //   in=0.556641 val=0.507927
    (addr==286) ? 8546601 :  //   in=0.558594 val=0.509417
    (addr==287) ? 8571555 :  //   in=0.560547 val=0.510905
    (addr==288) ? 8596468 :  //   in=0.562500 val=0.512389
    (addr==289) ? 8621339 :  //   in=0.564453 val=0.513872
    (addr==290) ? 8646169 :  //   in=0.566406 val=0.515352
    (addr==291) ? 8670957 :  //   in=0.568359 val=0.516829
    (addr==292) ? 8695704 :  //   in=0.570312 val=0.518304
    (addr==293) ? 8720409 :  //   in=0.572266 val=0.519777
    (addr==294) ? 8745072 :  //   in=0.574219 val=0.521247
    (addr==295) ? 8769694 :  //   in=0.576172 val=0.522715
    (addr==296) ? 8794274 :  //   in=0.578125 val=0.524180
    (addr==297) ? 8818813 :  //   in=0.580078 val=0.525642
    (addr==298) ? 8843310 :  //   in=0.582031 val=0.527102
    (addr==299) ? 8867766 :  //   in=0.583984 val=0.528560
    (addr==300) ? 8892180 :  //   in=0.585938 val=0.530015
    (addr==301) ? 8916552 :  //   in=0.587891 val=0.531468
    (addr==302) ? 8940883 :  //   in=0.589844 val=0.532918
    (addr==303) ? 8965173 :  //   in=0.591797 val=0.534366
    (addr==304) ? 8989420 :  //   in=0.593750 val=0.535811
    (addr==305) ? 9013627 :  //   in=0.595703 val=0.537254
    (addr==306) ? 9037791 :  //   in=0.597656 val=0.538694
    (addr==307) ? 9061915 :  //   in=0.599609 val=0.540132
    (addr==308) ? 9085996 :  //   in=0.601562 val=0.541568
    (addr==309) ? 9110036 :  //   in=0.603516 val=0.543001
    (addr==310) ? 9134035 :  //   in=0.605469 val=0.544431
    (addr==311) ? 9157992 :  //   in=0.607422 val=0.545859
    (addr==312) ? 9181908 :  //   in=0.609375 val=0.547284
    (addr==313) ? 9205782 :  //   in=0.611328 val=0.548707
    (addr==314) ? 9229615 :  //   in=0.613281 val=0.550128
    (addr==315) ? 9253406 :  //   in=0.615234 val=0.551546
    (addr==316) ? 9277156 :  //   in=0.617188 val=0.552962
    (addr==317) ? 9300864 :  //   in=0.619141 val=0.554375
    (addr==318) ? 9324531 :  //   in=0.621094 val=0.555785
    (addr==319) ? 9348157 :  //   in=0.623047 val=0.557194
    (addr==320) ? 9371741 :  //   in=0.625000 val=0.558599
    (addr==321) ? 9395284 :  //   in=0.626953 val=0.560003
    (addr==322) ? 9418785 :  //   in=0.628906 val=0.561403
    (addr==323) ? 9442245 :  //   in=0.630859 val=0.562802
    (addr==324) ? 9465664 :  //   in=0.632812 val=0.564198
    (addr==325) ? 9489042 :  //   in=0.634766 val=0.565591
    (addr==326) ? 9512378 :  //   in=0.636719 val=0.566982
    (addr==327) ? 9535673 :  //   in=0.638672 val=0.568370
    (addr==328) ? 9558927 :  //   in=0.640625 val=0.569756
    (addr==329) ? 9582139 :  //   in=0.642578 val=0.571140
    (addr==330) ? 9605310 :  //   in=0.644531 val=0.572521
    (addr==331) ? 9628441 :  //   in=0.646484 val=0.573900
    (addr==332) ? 9651530 :  //   in=0.648438 val=0.575276
    (addr==333) ? 9674577 :  //   in=0.650391 val=0.576650
    (addr==334) ? 9697584 :  //   in=0.652344 val=0.578021
    (addr==335) ? 9720550 :  //   in=0.654297 val=0.579390
    (addr==336) ? 9743474 :  //   in=0.656250 val=0.580756
    (addr==337) ? 9766358 :  //   in=0.658203 val=0.582120
    (addr==338) ? 9789200 :  //   in=0.660156 val=0.583482
    (addr==339) ? 9812002 :  //   in=0.662109 val=0.584841
    (addr==340) ? 9834762 :  //   in=0.664062 val=0.586198
    (addr==341) ? 9857482 :  //   in=0.666016 val=0.587552
    (addr==342) ? 9880161 :  //   in=0.667969 val=0.588904
    (addr==343) ? 9902799 :  //   in=0.669922 val=0.590253
    (addr==344) ? 9925396 :  //   in=0.671875 val=0.591600
    (addr==345) ? 9947952 :  //   in=0.673828 val=0.592944
    (addr==346) ? 9970467 :  //   in=0.675781 val=0.594286
    (addr==347) ? 9992942 :  //   in=0.677734 val=0.595626
    (addr==348) ? 10015376 :  //   in=0.679688 val=0.596963
    (addr==349) ? 10037769 :  //   in=0.681641 val=0.598298
    (addr==350) ? 10060121 :  //   in=0.683594 val=0.599630
    (addr==351) ? 10082433 :  //   in=0.685547 val=0.600960
    (addr==352) ? 10104704 :  //   in=0.687500 val=0.602287
    (addr==353) ? 10126935 :  //   in=0.689453 val=0.603612
    (addr==354) ? 10149125 :  //   in=0.691406 val=0.604935
    (addr==355) ? 10171275 :  //   in=0.693359 val=0.606255
    (addr==356) ? 10193384 :  //   in=0.695312 val=0.607573
    (addr==357) ? 10215453 :  //   in=0.697266 val=0.608888
    (addr==358) ? 10237481 :  //   in=0.699219 val=0.610201
    (addr==359) ? 10259469 :  //   in=0.701172 val=0.611512
    (addr==360) ? 10281416 :  //   in=0.703125 val=0.612820
    (addr==361) ? 10303324 :  //   in=0.705078 val=0.614126
    (addr==362) ? 10325191 :  //   in=0.707031 val=0.615429
    (addr==363) ? 10347017 :  //   in=0.708984 val=0.616730
    (addr==364) ? 10368804 :  //   in=0.710938 val=0.618029
    (addr==365) ? 10390550 :  //   in=0.712891 val=0.619325
    (addr==366) ? 10412257 :  //   in=0.714844 val=0.620619
    (addr==367) ? 10433923 :  //   in=0.716797 val=0.621910
    (addr==368) ? 10455549 :  //   in=0.718750 val=0.623199
    (addr==369) ? 10477135 :  //   in=0.720703 val=0.624486
    (addr==370) ? 10498682 :  //   in=0.722656 val=0.625770
    (addr==371) ? 10520188 :  //   in=0.724609 val=0.627052
    (addr==372) ? 10541655 :  //   in=0.726562 val=0.628332
    (addr==373) ? 10563081 :  //   in=0.728516 val=0.629609
    (addr==374) ? 10584468 :  //   in=0.730469 val=0.630883
    (addr==375) ? 10605815 :  //   in=0.732422 val=0.632156
    (addr==376) ? 10627122 :  //   in=0.734375 val=0.633426
    (addr==377) ? 10648390 :  //   in=0.736328 val=0.634694
    (addr==378) ? 10669618 :  //   in=0.738281 val=0.635959
    (addr==379) ? 10690807 :  //   in=0.740234 val=0.637222
    (addr==380) ? 10711955 :  //   in=0.742188 val=0.638482
    (addr==381) ? 10733065 :  //   in=0.744141 val=0.639741
    (addr==382) ? 10754135 :  //   in=0.746094 val=0.640996
    (addr==383) ? 10775165 :  //   in=0.748047 val=0.642250
    (addr==384) ? 10796157 :  //   in=0.750000 val=0.643501
    (addr==385) ? 10817108 :  //   in=0.751953 val=0.644750
    (addr==386) ? 10838021 :  //   in=0.753906 val=0.645996
    (addr==387) ? 10858894 :  //   in=0.755859 val=0.647241
    (addr==388) ? 10879729 :  //   in=0.757812 val=0.648482
    (addr==389) ? 10900524 :  //   in=0.759766 val=0.649722
    (addr==390) ? 10921280 :  //   in=0.761719 val=0.650959
    (addr==391) ? 10941996 :  //   in=0.763672 val=0.652194
    (addr==392) ? 10962674 :  //   in=0.765625 val=0.653426
    (addr==393) ? 10983313 :  //   in=0.767578 val=0.654657
    (addr==394) ? 11003913 :  //   in=0.769531 val=0.655884
    (addr==395) ? 11024475 :  //   in=0.771484 val=0.657110
    (addr==396) ? 11044997 :  //   in=0.773438 val=0.658333
    (addr==397) ? 11065481 :  //   in=0.775391 val=0.659554
    (addr==398) ? 11085925 :  //   in=0.777344 val=0.660773
    (addr==399) ? 11106332 :  //   in=0.779297 val=0.661989
    (addr==400) ? 11126699 :  //   in=0.781250 val=0.663203
    (addr==401) ? 11147028 :  //   in=0.783203 val=0.664415
    (addr==402) ? 11167319 :  //   in=0.785156 val=0.665624
    (addr==403) ? 11187571 :  //   in=0.787109 val=0.666831
    (addr==404) ? 11207785 :  //   in=0.789062 val=0.668036
    (addr==405) ? 11227960 :  //   in=0.791016 val=0.669239
    (addr==406) ? 11248097 :  //   in=0.792969 val=0.670439
    (addr==407) ? 11268196 :  //   in=0.794922 val=0.671637
    (addr==408) ? 11288256 :  //   in=0.796875 val=0.672833
    (addr==409) ? 11308279 :  //   in=0.798828 val=0.674026
    (addr==410) ? 11328263 :  //   in=0.800781 val=0.675217
    (addr==411) ? 11348209 :  //   in=0.802734 val=0.676406
    (addr==412) ? 11368118 :  //   in=0.804688 val=0.677593
    (addr==413) ? 11387988 :  //   in=0.806641 val=0.678777
    (addr==414) ? 11407820 :  //   in=0.808594 val=0.679959
    (addr==415) ? 11427615 :  //   in=0.810547 val=0.681139
    (addr==416) ? 11447372 :  //   in=0.812500 val=0.682317
    (addr==417) ? 11467091 :  //   in=0.814453 val=0.683492
    (addr==418) ? 11486772 :  //   in=0.816406 val=0.684665
    (addr==419) ? 11506416 :  //   in=0.818359 val=0.685836
    (addr==420) ? 11526022 :  //   in=0.820312 val=0.687004
    (addr==421) ? 11545591 :  //   in=0.822266 val=0.688171
    (addr==422) ? 11565122 :  //   in=0.824219 val=0.689335
    (addr==423) ? 11584616 :  //   in=0.826172 val=0.690497
    (addr==424) ? 11604072 :  //   in=0.828125 val=0.691657
    (addr==425) ? 11623491 :  //   in=0.830078 val=0.692814
    (addr==426) ? 11642873 :  //   in=0.832031 val=0.693969
    (addr==427) ? 11662218 :  //   in=0.833984 val=0.695122
    (addr==428) ? 11681525 :  //   in=0.835938 val=0.696273
    (addr==429) ? 11700796 :  //   in=0.837891 val=0.697422
    (addr==430) ? 11720029 :  //   in=0.839844 val=0.698568
    (addr==431) ? 11739226 :  //   in=0.841797 val=0.699712
    (addr==432) ? 11758385 :  //   in=0.843750 val=0.700854
    (addr==433) ? 11777508 :  //   in=0.845703 val=0.701994
    (addr==434) ? 11796594 :  //   in=0.847656 val=0.703132
    (addr==435) ? 11815643 :  //   in=0.849609 val=0.704267
    (addr==436) ? 11834656 :  //   in=0.851562 val=0.705400
    (addr==437) ? 11853632 :  //   in=0.853516 val=0.706532
    (addr==438) ? 11872571 :  //   in=0.855469 val=0.707660
    (addr==439) ? 11891474 :  //   in=0.857422 val=0.708787
    (addr==440) ? 11910340 :  //   in=0.859375 val=0.709912
    (addr==441) ? 11929170 :  //   in=0.861328 val=0.711034
    (addr==442) ? 11947964 :  //   in=0.863281 val=0.712154
    (addr==443) ? 11966721 :  //   in=0.865234 val=0.713272
    (addr==444) ? 11985442 :  //   in=0.867188 val=0.714388
    (addr==445) ? 12004127 :  //   in=0.869141 val=0.715502
    (addr==446) ? 12022776 :  //   in=0.871094 val=0.716613
    (addr==447) ? 12041389 :  //   in=0.873047 val=0.717723
    (addr==448) ? 12059966 :  //   in=0.875000 val=0.718830
    (addr==449) ? 12078507 :  //   in=0.876953 val=0.719935
    (addr==450) ? 12097012 :  //   in=0.878906 val=0.721038
    (addr==451) ? 12115481 :  //   in=0.880859 val=0.722139
    (addr==452) ? 12133914 :  //   in=0.882812 val=0.723238
    (addr==453) ? 12152312 :  //   in=0.884766 val=0.724334
    (addr==454) ? 12170674 :  //   in=0.886719 val=0.725429
    (addr==455) ? 12189001 :  //   in=0.888672 val=0.726521
    (addr==456) ? 12207292 :  //   in=0.890625 val=0.727611
    (addr==457) ? 12225548 :  //   in=0.892578 val=0.728699
    (addr==458) ? 12243768 :  //   in=0.894531 val=0.729785
    (addr==459) ? 12261953 :  //   in=0.896484 val=0.730869
    (addr==460) ? 12280102 :  //   in=0.898438 val=0.731951
    (addr==461) ? 12298217 :  //   in=0.900391 val=0.733031
    (addr==462) ? 12316296 :  //   in=0.902344 val=0.734108
    (addr==463) ? 12334340 :  //   in=0.904297 val=0.735184
    (addr==464) ? 12352349 :  //   in=0.906250 val=0.736257
    (addr==465) ? 12370324 :  //   in=0.908203 val=0.737329
    (addr==466) ? 12388263 :  //   in=0.910156 val=0.738398
    (addr==467) ? 12406167 :  //   in=0.912109 val=0.739465
    (addr==468) ? 12424037 :  //   in=0.914062 val=0.740530
    (addr==469) ? 12441872 :  //   in=0.916016 val=0.741593
    (addr==470) ? 12459672 :  //   in=0.917969 val=0.742654
    (addr==471) ? 12477438 :  //   in=0.919922 val=0.743713
    (addr==472) ? 12495169 :  //   in=0.921875 val=0.744770
    (addr==473) ? 12512865 :  //   in=0.923828 val=0.745825
    (addr==474) ? 12530528 :  //   in=0.925781 val=0.746878
    (addr==475) ? 12548155 :  //   in=0.927734 val=0.747928
    (addr==476) ? 12565749 :  //   in=0.929688 val=0.748977
    (addr==477) ? 12583308 :  //   in=0.931641 val=0.750024
    (addr==478) ? 12600833 :  //   in=0.933594 val=0.751068
    (addr==479) ? 12618324 :  //   in=0.935547 val=0.752111
    (addr==480) ? 12635781 :  //   in=0.937500 val=0.753151
    (addr==481) ? 12653204 :  //   in=0.939453 val=0.754190
    (addr==482) ? 12670593 :  //   in=0.941406 val=0.755226
    (addr==483) ? 12687948 :  //   in=0.943359 val=0.756261
    (addr==484) ? 12705270 :  //   in=0.945312 val=0.757293
    (addr==485) ? 12722557 :  //   in=0.947266 val=0.758324
    (addr==486) ? 12739811 :  //   in=0.949219 val=0.759352
    (addr==487) ? 12757031 :  //   in=0.951172 val=0.760378
    (addr==488) ? 12774218 :  //   in=0.953125 val=0.761403
    (addr==489) ? 12791371 :  //   in=0.955078 val=0.762425
    (addr==490) ? 12808491 :  //   in=0.957031 val=0.763446
    (addr==491) ? 12825578 :  //   in=0.958984 val=0.764464
    (addr==492) ? 12842631 :  //   in=0.960938 val=0.765480
    (addr==493) ? 12859651 :  //   in=0.962891 val=0.766495
    (addr==494) ? 12876637 :  //   in=0.964844 val=0.767507
    (addr==495) ? 12893591 :  //   in=0.966797 val=0.768518
    (addr==496) ? 12910511 :  //   in=0.968750 val=0.769526
    (addr==497) ? 12927399 :  //   in=0.970703 val=0.770533
    (addr==498) ? 12944254 :  //   in=0.972656 val=0.771538
    (addr==499) ? 12961075 :  //   in=0.974609 val=0.772540
    (addr==500) ? 12977864 :  //   in=0.976562 val=0.773541
    (addr==501) ? 12994620 :  //   in=0.978516 val=0.774540
    (addr==502) ? 13011344 :  //   in=0.980469 val=0.775537
    (addr==503) ? 13028035 :  //   in=0.982422 val=0.776531
    (addr==504) ? 13044693 :  //   in=0.984375 val=0.777524
    (addr==505) ? 13061319 :  //   in=0.986328 val=0.778515
    (addr==506) ? 13077912 :  //   in=0.988281 val=0.779504
    (addr==507) ? 13094473 :  //   in=0.990234 val=0.780491
    (addr==508) ? 13111001 :  //   in=0.992188 val=0.781477
    (addr==509) ? 13127498 :  //   in=0.994141 val=0.782460
    (addr==510) ? 13143962 :  //   in=0.996094 val=0.783441
    (addr==511) ? 13160394 :  //   in=0.998047 val=0.784421
    (addr==512) ? 13176794 :  //   in=1.000000 val=0.785398
    (addr==513) ? 13193162 :  //   in=1.001953 val=0.786374
    (addr==514) ? 13209498 :  //   in=1.003906 val=0.787347
    (addr==515) ? 13225802 :  //   in=1.005859 val=0.788319
    (addr==516) ? 13242075 :  //   in=1.007812 val=0.789289
    (addr==517) ? 13258315 :  //   in=1.009766 val=0.790257
    (addr==518) ? 13274524 :  //   in=1.011719 val=0.791223
    (addr==519) ? 13290702 :  //   in=1.013672 val=0.792188
    (addr==520) ? 13306847 :  //   in=1.015625 val=0.793150
    (addr==521) ? 13322962 :  //   in=1.017578 val=0.794110
    (addr==522) ? 13339045 :  //   in=1.019531 val=0.795069
    (addr==523) ? 13355096 :  //   in=1.021484 val=0.796026
    (addr==524) ? 13371116 :  //   in=1.023438 val=0.796981
    (addr==525) ? 13387105 :  //   in=1.025391 val=0.797934
    (addr==526) ? 13403063 :  //   in=1.027344 val=0.798885
    (addr==527) ? 13418989 :  //   in=1.029297 val=0.799834
    (addr==528) ? 13434885 :  //   in=1.031250 val=0.800782
    (addr==529) ? 13450749 :  //   in=1.033203 val=0.801727
    (addr==530) ? 13466583 :  //   in=1.035156 val=0.802671
    (addr==531) ? 13482386 :  //   in=1.037109 val=0.803613
    (addr==532) ? 13498157 :  //   in=1.039062 val=0.804553
    (addr==533) ? 13513899 :  //   in=1.041016 val=0.805491
    (addr==534) ? 13529609 :  //   in=1.042969 val=0.806428
    (addr==535) ? 13545289 :  //   in=1.044922 val=0.807362
    (addr==536) ? 13560938 :  //   in=1.046875 val=0.808295
    (addr==537) ? 13576557 :  //   in=1.048828 val=0.809226
    (addr==538) ? 13592145 :  //   in=1.050781 val=0.810155
    (addr==539) ? 13607703 :  //   in=1.052734 val=0.811082
    (addr==540) ? 13623231 :  //   in=1.054688 val=0.812008
    (addr==541) ? 13638728 :  //   in=1.056641 val=0.812932
    (addr==542) ? 13654195 :  //   in=1.058594 val=0.813853
    (addr==543) ? 13669632 :  //   in=1.060547 val=0.814774
    (addr==544) ? 13685039 :  //   in=1.062500 val=0.815692
    (addr==545) ? 13700416 :  //   in=1.064453 val=0.816608
    (addr==546) ? 13715763 :  //   in=1.066406 val=0.817523
    (addr==547) ? 13731080 :  //   in=1.068359 val=0.818436
    (addr==548) ? 13746367 :  //   in=1.070312 val=0.819347
    (addr==549) ? 13761625 :  //   in=1.072266 val=0.820257
    (addr==550) ? 13776853 :  //   in=1.074219 val=0.821164
    (addr==551) ? 13792051 :  //   in=1.076172 val=0.822070
    (addr==552) ? 13807220 :  //   in=1.078125 val=0.822974
    (addr==553) ? 13822359 :  //   in=1.080078 val=0.823877
    (addr==554) ? 13837468 :  //   in=1.082031 val=0.824777
    (addr==555) ? 13852549 :  //   in=1.083984 val=0.825676
    (addr==556) ? 13867600 :  //   in=1.085938 val=0.826573
    (addr==557) ? 13882621 :  //   in=1.087891 val=0.827469
    (addr==558) ? 13897614 :  //   in=1.089844 val=0.828362
    (addr==559) ? 13912577 :  //   in=1.091797 val=0.829254
    (addr==560) ? 13927511 :  //   in=1.093750 val=0.830144
    (addr==561) ? 13942417 :  //   in=1.095703 val=0.831033
    (addr==562) ? 13957293 :  //   in=1.097656 val=0.831920
    (addr==563) ? 13972140 :  //   in=1.099609 val=0.832804
    (addr==564) ? 13986959 :  //   in=1.101562 val=0.833688
    (addr==565) ? 14001748 :  //   in=1.103516 val=0.834569
    (addr==566) ? 14016509 :  //   in=1.105469 val=0.835449
    (addr==567) ? 14031242 :  //   in=1.107422 val=0.836327
    (addr==568) ? 14045945 :  //   in=1.109375 val=0.837204
    (addr==569) ? 14060621 :  //   in=1.111328 val=0.838078
    (addr==570) ? 14075267 :  //   in=1.113281 val=0.838951
    (addr==571) ? 14089886 :  //   in=1.115234 val=0.839823
    (addr==572) ? 14104476 :  //   in=1.117188 val=0.840692
    (addr==573) ? 14119037 :  //   in=1.119141 val=0.841560
    (addr==574) ? 14133571 :  //   in=1.121094 val=0.842426
    (addr==575) ? 14148076 :  //   in=1.123047 val=0.843291
    (addr==576) ? 14162553 :  //   in=1.125000 val=0.844154
    (addr==577) ? 14177002 :  //   in=1.126953 val=0.845015
    (addr==578) ? 14191423 :  //   in=1.128906 val=0.845875
    (addr==579) ? 14205817 :  //   in=1.130859 val=0.846733
    (addr==580) ? 14220182 :  //   in=1.132812 val=0.847589
    (addr==581) ? 14234519 :  //   in=1.134766 val=0.848444
    (addr==582) ? 14248829 :  //   in=1.136719 val=0.849296
    (addr==583) ? 14263111 :  //   in=1.138672 val=0.850148
    (addr==584) ? 14277366 :  //   in=1.140625 val=0.850997
    (addr==585) ? 14291592 :  //   in=1.142578 val=0.851845
    (addr==586) ? 14305792 :  //   in=1.144531 val=0.852692
    (addr==587) ? 14319964 :  //   in=1.146484 val=0.853536
    (addr==588) ? 14334108 :  //   in=1.148438 val=0.854379
    (addr==589) ? 14348225 :  //   in=1.150391 val=0.855221
    (addr==590) ? 14362315 :  //   in=1.152344 val=0.856061
    (addr==591) ? 14376378 :  //   in=1.154297 val=0.856899
    (addr==592) ? 14390413 :  //   in=1.156250 val=0.857735
    (addr==593) ? 14404422 :  //   in=1.158203 val=0.858570
    (addr==594) ? 14418403 :  //   in=1.160156 val=0.859404
    (addr==595) ? 14432357 :  //   in=1.162109 val=0.860236
    (addr==596) ? 14446285 :  //   in=1.164062 val=0.861066
    (addr==597) ? 14460185 :  //   in=1.166016 val=0.861894
    (addr==598) ? 14474059 :  //   in=1.167969 val=0.862721
    (addr==599) ? 14487906 :  //   in=1.169922 val=0.863547
    (addr==600) ? 14501726 :  //   in=1.171875 val=0.864370
    (addr==601) ? 14515520 :  //   in=1.173828 val=0.865192
    (addr==602) ? 14529287 :  //   in=1.175781 val=0.866013
    (addr==603) ? 14543028 :  //   in=1.177734 val=0.866832
    (addr==604) ? 14556742 :  //   in=1.179688 val=0.867649
    (addr==605) ? 14570430 :  //   in=1.181641 val=0.868465
    (addr==606) ? 14584091 :  //   in=1.183594 val=0.869280
    (addr==607) ? 14597726 :  //   in=1.185547 val=0.870092
    (addr==608) ? 14611335 :  //   in=1.187500 val=0.870903
    (addr==609) ? 14624918 :  //   in=1.189453 val=0.871713
    (addr==610) ? 14638474 :  //   in=1.191406 val=0.872521
    (addr==611) ? 14652005 :  //   in=1.193359 val=0.873328
    (addr==612) ? 14665509 :  //   in=1.195312 val=0.874133
    (addr==613) ? 14678988 :  //   in=1.197266 val=0.874936
    (addr==614) ? 14692441 :  //   in=1.199219 val=0.875738
    (addr==615) ? 14705868 :  //   in=1.201172 val=0.876538
    (addr==616) ? 14719269 :  //   in=1.203125 val=0.877337
    (addr==617) ? 14732644 :  //   in=1.205078 val=0.878134
    (addr==618) ? 14745994 :  //   in=1.207031 val=0.878930
    (addr==619) ? 14759318 :  //   in=1.208984 val=0.879724
    (addr==620) ? 14772617 :  //   in=1.210938 val=0.880517
    (addr==621) ? 14785890 :  //   in=1.212891 val=0.881308
    (addr==622) ? 14799138 :  //   in=1.214844 val=0.882097
    (addr==623) ? 14812360 :  //   in=1.216797 val=0.882886
    (addr==624) ? 14825557 :  //   in=1.218750 val=0.883672
    (addr==625) ? 14838729 :  //   in=1.220703 val=0.884457
    (addr==626) ? 14851876 :  //   in=1.222656 val=0.885241
    (addr==627) ? 14864997 :  //   in=1.224609 val=0.886023
    (addr==628) ? 14878094 :  //   in=1.226562 val=0.886804
    (addr==629) ? 14891165 :  //   in=1.228516 val=0.887583
    (addr==630) ? 14904212 :  //   in=1.230469 val=0.888360
    (addr==631) ? 14917233 :  //   in=1.232422 val=0.889136
    (addr==632) ? 14930230 :  //   in=1.234375 val=0.889911
    (addr==633) ? 14943202 :  //   in=1.236328 val=0.890684
    (addr==634) ? 14956149 :  //   in=1.238281 val=0.891456
    (addr==635) ? 14969071 :  //   in=1.240234 val=0.892226
    (addr==636) ? 14981969 :  //   in=1.242188 val=0.892995
    (addr==637) ? 14994842 :  //   in=1.244141 val=0.893762
    (addr==638) ? 15007690 :  //   in=1.246094 val=0.894528
    (addr==639) ? 15020515 :  //   in=1.248047 val=0.895292
    (addr==640) ? 15033314 :  //   in=1.250000 val=0.896055
    (addr==641) ? 15046090 :  //   in=1.251953 val=0.896817
    (addr==642) ? 15058841 :  //   in=1.253906 val=0.897577
    (addr==643) ? 15071567 :  //   in=1.255859 val=0.898335
    (addr==644) ? 15084270 :  //   in=1.257812 val=0.899093
    (addr==645) ? 15096948 :  //   in=1.259766 val=0.899848
    (addr==646) ? 15109603 :  //   in=1.261719 val=0.900603
    (addr==647) ? 15122233 :  //   in=1.263672 val=0.901355
    (addr==648) ? 15134839 :  //   in=1.265625 val=0.902107
    (addr==649) ? 15147422 :  //   in=1.267578 val=0.902857
    (addr==650) ? 15159980 :  //   in=1.269531 val=0.903605
    (addr==651) ? 15172515 :  //   in=1.271484 val=0.904352
    (addr==652) ? 15185026 :  //   in=1.273438 val=0.905098
    (addr==653) ? 15197513 :  //   in=1.275391 val=0.905842
    (addr==654) ? 15209976 :  //   in=1.277344 val=0.906585
    (addr==655) ? 15222416 :  //   in=1.279297 val=0.907327
    (addr==656) ? 15234833 :  //   in=1.281250 val=0.908067
    (addr==657) ? 15247226 :  //   in=1.283203 val=0.908805
    (addr==658) ? 15259595 :  //   in=1.285156 val=0.909543
    (addr==659) ? 15271941 :  //   in=1.287109 val=0.910279
    (addr==660) ? 15284264 :  //   in=1.289062 val=0.911013
    (addr==661) ? 15296563 :  //   in=1.291016 val=0.911746
    (addr==662) ? 15308839 :  //   in=1.292969 val=0.912478
    (addr==663) ? 15321092 :  //   in=1.294922 val=0.913208
    (addr==664) ? 15333322 :  //   in=1.296875 val=0.913937
    (addr==665) ? 15345529 :  //   in=1.298828 val=0.914665
    (addr==666) ? 15357712 :  //   in=1.300781 val=0.915391
    (addr==667) ? 15369873 :  //   in=1.302734 val=0.916116
    (addr==668) ? 15382011 :  //   in=1.304688 val=0.916839
    (addr==669) ? 15394126 :  //   in=1.306641 val=0.917561
    (addr==670) ? 15406218 :  //   in=1.308594 val=0.918282
    (addr==671) ? 15418287 :  //   in=1.310547 val=0.919002
    (addr==672) ? 15430334 :  //   in=1.312500 val=0.919720
    (addr==673) ? 15442358 :  //   in=1.314453 val=0.920436
    (addr==674) ? 15454359 :  //   in=1.316406 val=0.921152
    (addr==675) ? 15466338 :  //   in=1.318359 val=0.921866
    (addr==676) ? 15478294 :  //   in=1.320312 val=0.922578
    (addr==677) ? 15490228 :  //   in=1.322266 val=0.923290
    (addr==678) ? 15502140 :  //   in=1.324219 val=0.924000
    (addr==679) ? 15514029 :  //   in=1.326172 val=0.924708
    (addr==680) ? 15525896 :  //   in=1.328125 val=0.925416
    (addr==681) ? 15537740 :  //   in=1.330078 val=0.926122
    (addr==682) ? 15549562 :  //   in=1.332031 val=0.926826
    (addr==683) ? 15561363 :  //   in=1.333984 val=0.927530
    (addr==684) ? 15573141 :  //   in=1.335938 val=0.928232
    (addr==685) ? 15584897 :  //   in=1.337891 val=0.928932
    (addr==686) ? 15596631 :  //   in=1.339844 val=0.929632
    (addr==687) ? 15608343 :  //   in=1.341797 val=0.930330
    (addr==688) ? 15620033 :  //   in=1.343750 val=0.931027
    (addr==689) ? 15631701 :  //   in=1.345703 val=0.931722
    (addr==690) ? 15643348 :  //   in=1.347656 val=0.932416
    (addr==691) ? 15654973 :  //   in=1.349609 val=0.933109
    (addr==692) ? 15666576 :  //   in=1.351562 val=0.933801
    (addr==693) ? 15678157 :  //   in=1.353516 val=0.934491
    (addr==694) ? 15689717 :  //   in=1.355469 val=0.935180
    (addr==695) ? 15701255 :  //   in=1.357422 val=0.935868
    (addr==696) ? 15712772 :  //   in=1.359375 val=0.936554
    (addr==697) ? 15724267 :  //   in=1.361328 val=0.937239
    (addr==698) ? 15735741 :  //   in=1.363281 val=0.937923
    (addr==699) ? 15747194 :  //   in=1.365234 val=0.938606
    (addr==700) ? 15758625 :  //   in=1.367188 val=0.939287
    (addr==701) ? 15770035 :  //   in=1.369141 val=0.939967
    (addr==702) ? 15781424 :  //   in=1.371094 val=0.940646
    (addr==703) ? 15792791 :  //   in=1.373047 val=0.941324
    (addr==704) ? 15804138 :  //   in=1.375000 val=0.942000
    (addr==705) ? 15815463 :  //   in=1.376953 val=0.942675
    (addr==706) ? 15826768 :  //   in=1.378906 val=0.943349
    (addr==707) ? 15838051 :  //   in=1.380859 val=0.944021
    (addr==708) ? 15849313 :  //   in=1.382812 val=0.944693
    (addr==709) ? 15860555 :  //   in=1.384766 val=0.945363
    (addr==710) ? 15871776 :  //   in=1.386719 val=0.946032
    (addr==711) ? 15882976 :  //   in=1.388672 val=0.946699
    (addr==712) ? 15894155 :  //   in=1.390625 val=0.947366
    (addr==713) ? 15905314 :  //   in=1.392578 val=0.948031
    (addr==714) ? 15916452 :  //   in=1.394531 val=0.948695
    (addr==715) ? 15927570 :  //   in=1.396484 val=0.949357
    (addr==716) ? 15938666 :  //   in=1.398438 val=0.950019
    (addr==717) ? 15949743 :  //   in=1.400391 val=0.950679
    (addr==718) ? 15960799 :  //   in=1.402344 val=0.951338
    (addr==719) ? 15971834 :  //   in=1.404297 val=0.951996
    (addr==720) ? 15982850 :  //   in=1.406250 val=0.952652
    (addr==721) ? 15993844 :  //   in=1.408203 val=0.953307
    (addr==722) ? 16004819 :  //   in=1.410156 val=0.953962
    (addr==723) ? 16015774 :  //   in=1.412109 val=0.954615
    (addr==724) ? 16026708 :  //   in=1.414062 val=0.955266
    (addr==725) ? 16037622 :  //   in=1.416016 val=0.955917
    (addr==726) ? 16048516 :  //   in=1.417969 val=0.956566
    (addr==727) ? 16059390 :  //   in=1.419922 val=0.957214
    (addr==728) ? 16070244 :  //   in=1.421875 val=0.957861
    (addr==729) ? 16081079 :  //   in=1.423828 val=0.958507
    (addr==730) ? 16091893 :  //   in=1.425781 val=0.959152
    (addr==731) ? 16102687 :  //   in=1.427734 val=0.959795
    (addr==732) ? 16113462 :  //   in=1.429688 val=0.960437
    (addr==733) ? 16124217 :  //   in=1.431641 val=0.961078
    (addr==734) ? 16134952 :  //   in=1.433594 val=0.961718
    (addr==735) ? 16145667 :  //   in=1.435547 val=0.962357
    (addr==736) ? 16156363 :  //   in=1.437500 val=0.962994
    (addr==737) ? 16167040 :  //   in=1.439453 val=0.963631
    (addr==738) ? 16177697 :  //   in=1.441406 val=0.964266
    (addr==739) ? 16188334 :  //   in=1.443359 val=0.964900
    (addr==740) ? 16198952 :  //   in=1.445312 val=0.965533
    (addr==741) ? 16209550 :  //   in=1.447266 val=0.966165
    (addr==742) ? 16220130 :  //   in=1.449219 val=0.966795
    (addr==743) ? 16230689 :  //   in=1.451172 val=0.967425
    (addr==744) ? 16241230 :  //   in=1.453125 val=0.968053
    (addr==745) ? 16251751 :  //   in=1.455078 val=0.968680
    (addr==746) ? 16262254 :  //   in=1.457031 val=0.969306
    (addr==747) ? 16272737 :  //   in=1.458984 val=0.969931
    (addr==748) ? 16283201 :  //   in=1.460938 val=0.970554
    (addr==749) ? 16293646 :  //   in=1.462891 val=0.971177
    (addr==750) ? 16304072 :  //   in=1.464844 val=0.971798
    (addr==751) ? 16314479 :  //   in=1.466797 val=0.972419
    (addr==752) ? 16324867 :  //   in=1.468750 val=0.973038
    (addr==753) ? 16335236 :  //   in=1.470703 val=0.973656
    (addr==754) ? 16345587 :  //   in=1.472656 val=0.974273
    (addr==755) ? 16355919 :  //   in=1.474609 val=0.974889
    (addr==756) ? 16366232 :  //   in=1.476562 val=0.975503
    (addr==757) ? 16376526 :  //   in=1.478516 val=0.976117
    (addr==758) ? 16386802 :  //   in=1.480469 val=0.976730
    (addr==759) ? 16397059 :  //   in=1.482422 val=0.977341
    (addr==760) ? 16407297 :  //   in=1.484375 val=0.977951
    (addr==761) ? 16417517 :  //   in=1.486328 val=0.978560
    (addr==762) ? 16427719 :  //   in=1.488281 val=0.979168
    (addr==763) ? 16437902 :  //   in=1.490234 val=0.979775
    (addr==764) ? 16448066 :  //   in=1.492188 val=0.980381
    (addr==765) ? 16458213 :  //   in=1.494141 val=0.980986
    (addr==766) ? 16468341 :  //   in=1.496094 val=0.981590
    (addr==767) ? 16478451 :  //   in=1.498047 val=0.982192
    (addr==768) ? 16488542 :  //   in=1.500000 val=0.982794
    (addr==769) ? 16498615 :  //   in=1.501953 val=0.983394
    (addr==770) ? 16508671 :  //   in=1.503906 val=0.983993
    (addr==771) ? 16518708 :  //   in=1.505859 val=0.984592
    (addr==772) ? 16528727 :  //   in=1.507812 val=0.985189
    (addr==773) ? 16538728 :  //   in=1.509766 val=0.985785
    (addr==774) ? 16548711 :  //   in=1.511719 val=0.986380
    (addr==775) ? 16558676 :  //   in=1.513672 val=0.986974
    (addr==776) ? 16568624 :  //   in=1.515625 val=0.987567
    (addr==777) ? 16578553 :  //   in=1.517578 val=0.988159
    (addr==778) ? 16588465 :  //   in=1.519531 val=0.988750
    (addr==779) ? 16598359 :  //   in=1.521484 val=0.989339
    (addr==780) ? 16608235 :  //   in=1.523438 val=0.989928
    (addr==781) ? 16618093 :  //   in=1.525391 val=0.990516
    (addr==782) ? 16627934 :  //   in=1.527344 val=0.991102
    (addr==783) ? 16637757 :  //   in=1.529297 val=0.991688
    (addr==784) ? 16647563 :  //   in=1.531250 val=0.992272
    (addr==785) ? 16657351 :  //   in=1.533203 val=0.992856
    (addr==786) ? 16667122 :  //   in=1.535156 val=0.993438
    (addr==787) ? 16676875 :  //   in=1.537109 val=0.994019
    (addr==788) ? 16686611 :  //   in=1.539062 val=0.994600
    (addr==789) ? 16696329 :  //   in=1.541016 val=0.995179
    (addr==790) ? 16706031 :  //   in=1.542969 val=0.995757
    (addr==791) ? 16715715 :  //   in=1.544922 val=0.996334
    (addr==792) ? 16725381 :  //   in=1.546875 val=0.996910
    (addr==793) ? 16735031 :  //   in=1.548828 val=0.997486
    (addr==794) ? 16744663 :  //   in=1.550781 val=0.998060
    (addr==795) ? 16754278 :  //   in=1.552734 val=0.998633
    (addr==796) ? 16763876 :  //   in=1.554688 val=0.999205
    (addr==797) ? 16773457 :  //   in=1.556641 val=0.999776
    (addr==798) ? 16783021 :  //   in=1.558594 val=1.000346
    (addr==799) ? 16792568 :  //   in=1.560547 val=1.000915
    (addr==800) ? 16802098 :  //   in=1.562500 val=1.001483
    (addr==801) ? 16811612 :  //   in=1.564453 val=1.002050
    (addr==802) ? 16821108 :  //   in=1.566406 val=1.002616
    (addr==803) ? 16830588 :  //   in=1.568359 val=1.003181
    (addr==804) ? 16840050 :  //   in=1.570312 val=1.003745
    (addr==805) ? 16849497 :  //   in=1.572266 val=1.004308
    (addr==806) ? 16858926 :  //   in=1.574219 val=1.004870
    (addr==807) ? 16868339 :  //   in=1.576172 val=1.005431
    (addr==808) ? 16877735 :  //   in=1.578125 val=1.005991
    (addr==809) ? 16887114 :  //   in=1.580078 val=1.006550
    (addr==810) ? 16896477 :  //   in=1.582031 val=1.007109
    (addr==811) ? 16905824 :  //   in=1.583984 val=1.007666
    (addr==812) ? 16915154 :  //   in=1.585938 val=1.008222
    (addr==813) ? 16924467 :  //   in=1.587891 val=1.008777
    (addr==814) ? 16933765 :  //   in=1.589844 val=1.009331
    (addr==815) ? 16943046 :  //   in=1.591797 val=1.009884
    (addr==816) ? 16952310 :  //   in=1.593750 val=1.010436
    (addr==817) ? 16961558 :  //   in=1.595703 val=1.010988
    (addr==818) ? 16970790 :  //   in=1.597656 val=1.011538
    (addr==819) ? 16980006 :  //   in=1.599609 val=1.012087
    (addr==820) ? 16989206 :  //   in=1.601562 val=1.012636
    (addr==821) ? 16998389 :  //   in=1.603516 val=1.013183
    (addr==822) ? 17007557 :  //   in=1.605469 val=1.013729
    (addr==823) ? 17016708 :  //   in=1.607422 val=1.014275
    (addr==824) ? 17025843 :  //   in=1.609375 val=1.014819
    (addr==825) ? 17034963 :  //   in=1.611328 val=1.015363
    (addr==826) ? 17044066 :  //   in=1.613281 val=1.015906
    (addr==827) ? 17053154 :  //   in=1.615234 val=1.016447
    (addr==828) ? 17062225 :  //   in=1.617188 val=1.016988
    (addr==829) ? 17071281 :  //   in=1.619141 val=1.017528
    (addr==830) ? 17080321 :  //   in=1.621094 val=1.018067
    (addr==831) ? 17089345 :  //   in=1.623047 val=1.018604
    (addr==832) ? 17098354 :  //   in=1.625000 val=1.019141
    (addr==833) ? 17107347 :  //   in=1.626953 val=1.019677
    (addr==834) ? 17116324 :  //   in=1.628906 val=1.020212
    (addr==835) ? 17125285 :  //   in=1.630859 val=1.020747
    (addr==836) ? 17134231 :  //   in=1.632812 val=1.021280
    (addr==837) ? 17143162 :  //   in=1.634766 val=1.021812
    (addr==838) ? 17152077 :  //   in=1.636719 val=1.022343
    (addr==839) ? 17160976 :  //   in=1.638672 val=1.022874
    (addr==840) ? 17169860 :  //   in=1.640625 val=1.023403
    (addr==841) ? 17178729 :  //   in=1.642578 val=1.023932
    (addr==842) ? 17187582 :  //   in=1.644531 val=1.024460
    (addr==843) ? 17196420 :  //   in=1.646484 val=1.024987
    (addr==844) ? 17205242 :  //   in=1.648438 val=1.025512
    (addr==845) ? 17214049 :  //   in=1.650391 val=1.026037
    (addr==846) ? 17222841 :  //   in=1.652344 val=1.026561
    (addr==847) ? 17231618 :  //   in=1.654297 val=1.027085
    (addr==848) ? 17240380 :  //   in=1.656250 val=1.027607
    (addr==849) ? 17249126 :  //   in=1.658203 val=1.028128
    (addr==850) ? 17257858 :  //   in=1.660156 val=1.028649
    (addr==851) ? 17266574 :  //   in=1.662109 val=1.029168
    (addr==852) ? 17275276 :  //   in=1.664062 val=1.029687
    (addr==853) ? 17283962 :  //   in=1.666016 val=1.030204
    (addr==854) ? 17292633 :  //   in=1.667969 val=1.030721
    (addr==855) ? 17301290 :  //   in=1.669922 val=1.031237
    (addr==856) ? 17309931 :  //   in=1.671875 val=1.031752
    (addr==857) ? 17318558 :  //   in=1.673828 val=1.032267
    (addr==858) ? 17327170 :  //   in=1.675781 val=1.032780
    (addr==859) ? 17335767 :  //   in=1.677734 val=1.033292
    (addr==860) ? 17344349 :  //   in=1.679688 val=1.033804
    (addr==861) ? 17352917 :  //   in=1.681641 val=1.034314
    (addr==862) ? 17361470 :  //   in=1.683594 val=1.034824
    (addr==863) ? 17370008 :  //   in=1.685547 val=1.035333
    (addr==864) ? 17378532 :  //   in=1.687500 val=1.035841
    (addr==865) ? 17387041 :  //   in=1.689453 val=1.036348
    (addr==866) ? 17395536 :  //   in=1.691406 val=1.036855
    (addr==867) ? 17404015 :  //   in=1.693359 val=1.037360
    (addr==868) ? 17412481 :  //   in=1.695312 val=1.037865
    (addr==869) ? 17420932 :  //   in=1.697266 val=1.038368
    (addr==870) ? 17429369 :  //   in=1.699219 val=1.038871
    (addr==871) ? 17437791 :  //   in=1.701172 val=1.039373
    (addr==872) ? 17446199 :  //   in=1.703125 val=1.039875
    (addr==873) ? 17454592 :  //   in=1.705078 val=1.040375
    (addr==874) ? 17462971 :  //   in=1.707031 val=1.040874
    (addr==875) ? 17471336 :  //   in=1.708984 val=1.041373
    (addr==876) ? 17479687 :  //   in=1.710938 val=1.041871
    (addr==877) ? 17488024 :  //   in=1.712891 val=1.042367
    (addr==878) ? 17496346 :  //   in=1.714844 val=1.042864
    (addr==879) ? 17504654 :  //   in=1.716797 val=1.043359
    (addr==880) ? 17512948 :  //   in=1.718750 val=1.043853
    (addr==881) ? 17521228 :  //   in=1.720703 val=1.044347
    (addr==882) ? 17529495 :  //   in=1.722656 val=1.044839
    (addr==883) ? 17537747 :  //   in=1.724609 val=1.045331
    (addr==884) ? 17545985 :  //   in=1.726562 val=1.045822
    (addr==885) ? 17554209 :  //   in=1.728516 val=1.046312
    (addr==886) ? 17562419 :  //   in=1.730469 val=1.046802
    (addr==887) ? 17570615 :  //   in=1.732422 val=1.047290
    (addr==888) ? 17578798 :  //   in=1.734375 val=1.047778
    (addr==889) ? 17586966 :  //   in=1.736328 val=1.048265
    (addr==890) ? 17595121 :  //   in=1.738281 val=1.048751
    (addr==891) ? 17603262 :  //   in=1.740234 val=1.049236
    (addr==892) ? 17611389 :  //   in=1.742188 val=1.049721
    (addr==893) ? 17619503 :  //   in=1.744141 val=1.050204
    (addr==894) ? 17627603 :  //   in=1.746094 val=1.050687
    (addr==895) ? 17635690 :  //   in=1.748047 val=1.051169
    (addr==896) ? 17643762 :  //   in=1.750000 val=1.051650
    (addr==897) ? 17651821 :  //   in=1.751953 val=1.052131
    (addr==898) ? 17659867 :  //   in=1.753906 val=1.052610
    (addr==899) ? 17667899 :  //   in=1.755859 val=1.053089
    (addr==900) ? 17675918 :  //   in=1.757812 val=1.053567
    (addr==901) ? 17683923 :  //   in=1.759766 val=1.054044
    (addr==902) ? 17691915 :  //   in=1.761719 val=1.054520
    (addr==903) ? 17699893 :  //   in=1.763672 val=1.054996
    (addr==904) ? 17707858 :  //   in=1.765625 val=1.055471
    (addr==905) ? 17715810 :  //   in=1.767578 val=1.055945
    (addr==906) ? 17723748 :  //   in=1.769531 val=1.056418
    (addr==907) ? 17731674 :  //   in=1.771484 val=1.056890
    (addr==908) ? 17739585 :  //   in=1.773438 val=1.057362
    (addr==909) ? 17747484 :  //   in=1.775391 val=1.057833
    (addr==910) ? 17755370 :  //   in=1.777344 val=1.058303
    (addr==911) ? 17763242 :  //   in=1.779297 val=1.058772
    (addr==912) ? 17771101 :  //   in=1.781250 val=1.059240
    (addr==913) ? 17778947 :  //   in=1.783203 val=1.059708
    (addr==914) ? 17786780 :  //   in=1.785156 val=1.060175
    (addr==915) ? 17794600 :  //   in=1.787109 val=1.060641
    (addr==916) ? 17802407 :  //   in=1.789062 val=1.061106
    (addr==917) ? 17810201 :  //   in=1.791016 val=1.061571
    (addr==918) ? 17817982 :  //   in=1.792969 val=1.062035
    (addr==919) ? 17825751 :  //   in=1.794922 val=1.062498
    (addr==920) ? 17833506 :  //   in=1.796875 val=1.062960
    (addr==921) ? 17841248 :  //   in=1.798828 val=1.063421
    (addr==922) ? 17848978 :  //   in=1.800781 val=1.063882
    (addr==923) ? 17856695 :  //   in=1.802734 val=1.064342
    (addr==924) ? 17864399 :  //   in=1.804688 val=1.064801
    (addr==925) ? 17872090 :  //   in=1.806641 val=1.065260
    (addr==926) ? 17879768 :  //   in=1.808594 val=1.065717
    (addr==927) ? 17887434 :  //   in=1.810547 val=1.066174
    (addr==928) ? 17895088 :  //   in=1.812500 val=1.066630
    (addr==929) ? 17902728 :  //   in=1.814453 val=1.067086
    (addr==930) ? 17910356 :  //   in=1.816406 val=1.067540
    (addr==931) ? 17917971 :  //   in=1.818359 val=1.067994
    (addr==932) ? 17925574 :  //   in=1.820312 val=1.068448
    (addr==933) ? 17933164 :  //   in=1.822266 val=1.068900
    (addr==934) ? 17940742 :  //   in=1.824219 val=1.069352
    (addr==935) ? 17948308 :  //   in=1.826172 val=1.069803
    (addr==936) ? 17955861 :  //   in=1.828125 val=1.070253
    (addr==937) ? 17963401 :  //   in=1.830078 val=1.070702
    (addr==938) ? 17970929 :  //   in=1.832031 val=1.071151
    (addr==939) ? 17978445 :  //   in=1.833984 val=1.071599
    (addr==940) ? 17985948 :  //   in=1.835938 val=1.072046
    (addr==941) ? 17993439 :  //   in=1.837891 val=1.072493
    (addr==942) ? 18000918 :  //   in=1.839844 val=1.072938
    (addr==943) ? 18008385 :  //   in=1.841797 val=1.073383
    (addr==944) ? 18015839 :  //   in=1.843750 val=1.073828
    (addr==945) ? 18023281 :  //   in=1.845703 val=1.074271
    (addr==946) ? 18030711 :  //   in=1.847656 val=1.074714
    (addr==947) ? 18038129 :  //   in=1.849609 val=1.075156
    (addr==948) ? 18045535 :  //   in=1.851562 val=1.075598
    (addr==949) ? 18052929 :  //   in=1.853516 val=1.076038
    (addr==950) ? 18060310 :  //   in=1.855469 val=1.076478
    (addr==951) ? 18067680 :  //   in=1.857422 val=1.076918
    (addr==952) ? 18075037 :  //   in=1.859375 val=1.077356
    (addr==953) ? 18082383 :  //   in=1.861328 val=1.077794
    (addr==954) ? 18089717 :  //   in=1.863281 val=1.078231
    (addr==955) ? 18097038 :  //   in=1.865234 val=1.078668
    (addr==956) ? 18104348 :  //   in=1.867188 val=1.079103
    (addr==957) ? 18111646 :  //   in=1.869141 val=1.079538
    (addr==958) ? 18118932 :  //   in=1.871094 val=1.079973
    (addr==959) ? 18126206 :  //   in=1.873047 val=1.080406
    (addr==960) ? 18133469 :  //   in=1.875000 val=1.080839
    (addr==961) ? 18140720 :  //   in=1.876953 val=1.081271
    (addr==962) ? 18147959 :  //   in=1.878906 val=1.081703
    (addr==963) ? 18155186 :  //   in=1.880859 val=1.082133
    (addr==964) ? 18162401 :  //   in=1.882812 val=1.082564
    (addr==965) ? 18169605 :  //   in=1.884766 val=1.082993
    (addr==966) ? 18176797 :  //   in=1.886719 val=1.083422
    (addr==967) ? 18183978 :  //   in=1.888672 val=1.083850
    (addr==968) ? 18191147 :  //   in=1.890625 val=1.084277
    (addr==969) ? 18198305 :  //   in=1.892578 val=1.084704
    (addr==970) ? 18205450 :  //   in=1.894531 val=1.085129
    (addr==971) ? 18212585 :  //   in=1.896484 val=1.085555
    (addr==972) ? 18219708 :  //   in=1.898438 val=1.085979
    (addr==973) ? 18226819 :  //   in=1.900391 val=1.086403
    (addr==974) ? 18233919 :  //   in=1.902344 val=1.086826
    (addr==975) ? 18241008 :  //   in=1.904297 val=1.087249
    (addr==976) ? 18248085 :  //   in=1.906250 val=1.087671
    (addr==977) ? 18255151 :  //   in=1.908203 val=1.088092
    (addr==978) ? 18262206 :  //   in=1.910156 val=1.088512
    (addr==979) ? 18269249 :  //   in=1.912109 val=1.088932
    (addr==980) ? 18276281 :  //   in=1.914062 val=1.089351
    (addr==981) ? 18283301 :  //   in=1.916016 val=1.089770
    (addr==982) ? 18290311 :  //   in=1.917969 val=1.090188
    (addr==983) ? 18297309 :  //   in=1.919922 val=1.090605
    (addr==984) ? 18304296 :  //   in=1.921875 val=1.091021
    (addr==985) ? 18311272 :  //   in=1.923828 val=1.091437
    (addr==986) ? 18318236 :  //   in=1.925781 val=1.091852
    (addr==987) ? 18325190 :  //   in=1.927734 val=1.092266
    (addr==988) ? 18332132 :  //   in=1.929688 val=1.092680
    (addr==989) ? 18339064 :  //   in=1.931641 val=1.093093
    (addr==990) ? 18345984 :  //   in=1.933594 val=1.093506
    (addr==991) ? 18352894 :  //   in=1.935547 val=1.093918
    (addr==992) ? 18359792 :  //   in=1.937500 val=1.094329
    (addr==993) ? 18366679 :  //   in=1.939453 val=1.094739
    (addr==994) ? 18373556 :  //   in=1.941406 val=1.095149
    (addr==995) ? 18380421 :  //   in=1.943359 val=1.095559
    (addr==996) ? 18387276 :  //   in=1.945312 val=1.095967
    (addr==997) ? 18394120 :  //   in=1.947266 val=1.096375
    (addr==998) ? 18400952 :  //   in=1.949219 val=1.096782
    (addr==999) ? 18407774 :  //   in=1.951172 val=1.097189
    (addr==1000) ? 18414586 :  //   in=1.953125 val=1.097595
    (addr==1001) ? 18421386 :  //   in=1.955078 val=1.098000
    (addr==1002) ? 18428176 :  //   in=1.957031 val=1.098405
    (addr==1003) ? 18434955 :  //   in=1.958984 val=1.098809
    (addr==1004) ? 18441723 :  //   in=1.960938 val=1.099212
    (addr==1005) ? 18448481 :  //   in=1.962891 val=1.099615
    (addr==1006) ? 18455227 :  //   in=1.964844 val=1.100017
    (addr==1007) ? 18461964 :  //   in=1.966797 val=1.100419
    (addr==1008) ? 18468689 :  //   in=1.968750 val=1.100820
    (addr==1009) ? 18475404 :  //   in=1.970703 val=1.101220
    (addr==1010) ? 18482109 :  //   in=1.972656 val=1.101620
    (addr==1011) ? 18488802 :  //   in=1.974609 val=1.102019
    (addr==1012) ? 18495486 :  //   in=1.976562 val=1.102417
    (addr==1013) ? 18502159 :  //   in=1.978516 val=1.102815
    (addr==1014) ? 18508821 :  //   in=1.980469 val=1.103212
    (addr==1015) ? 18515473 :  //   in=1.982422 val=1.103608
    (addr==1016) ? 18522114 :  //   in=1.984375 val=1.104004
    (addr==1017) ? 18528745 :  //   in=1.986328 val=1.104399
    (addr==1018) ? 18535366 :  //   in=1.988281 val=1.104794
    (addr==1019) ? 18541976 :  //   in=1.990234 val=1.105188
    (addr==1020) ? 18548576 :  //   in=1.992188 val=1.105581
    (addr==1021) ? 18555166 :  //   in=1.994141 val=1.105974
    (addr==1022) ? 18561745 :  //   in=1.996094 val=1.106366
    (addr==1023) ? 18568314 :  //   in=1.998047 val=1.106758
25'bx;
assign lastone = 18574873;
endmodule
