
`timescale 1ns/1ps
module tb;
parameter IDWID=4; parameter DWID=64; parameter EXTRAS=8; parameter WSTRB=DWID/8;

integer    cycles;   initial cycles=0;
integer    errors;   initial errors=0;
integer    wrongs;   initial wrongs=0;
integer    Panics;   initial Panics=0;
integer    corrects; initial corrects=0;
reg [31:0] marker;   initial marker=0;
reg [31:0] marker0;   initial marker0=0;
reg [31:0] marker1;   initial marker1=0;
reg [31:0] marker2;   initial marker2=0;
reg [31:0] marker3;   initial marker3=0;
reg [31:0] Index;   initial Index=0;
integer    rqueuelen;   initial rqueuelen=0;
reg [31:0] seqptr;   initial seqptr=0;
reg [31:0] slv0_marker3;   initial slv0_marker3=0;
reg [31:0] slv1_marker3;   initial slv1_marker3=0;
reg [31:0] slv2_marker3;   initial slv2_marker3=0;
reg [31:0] slv3_marker3;   initial slv3_marker3=0;



reg clk; reg rst_n;
integer clk_HALFPERIOD = 100;
always begin
    clk = 0;
    #(clk_HALFPERIOD);
    clk = 1;
    #3;
    $python("negedge()");
    #3;
    $python("auxs()");
    #(clk_HALFPERIOD-6);
end
initial begin
    $dumpvars(0,tb);
    rst_n = 0;
    #100;
    rst_n = 1;
end

// reg  [2:0] slv0_awsize ; initial slv0_awsize = 0;
// reg  [2:0] slv0_arsize ; initial slv0_arsize = 0;

wire  [IDWID-1:0] slv0_arid ;
wire  [31:0] slv0_araddr ;
wire  [7:0] slv0_arlen ;
wire  [2:0] slv0_arsize ;
wire  [EXTRAS-1:0] slv0_arextras ;
wire  [1:0] slv0_arburst ;
wire  slv0_arvalid ;
reg  slv0_arready ;
reg  [IDWID-1:0] slv0_rid ;
reg  [DWID-1:0] slv0_rdata ;
reg  [1:0] slv0_rresp ;
reg  slv0_rlast ;
reg  slv0_rvalid ;
wire  slv0_rready ;

wire  [IDWID-1:0] slv0_awid ;
wire  [31:0] slv0_awaddr ;
wire  [7:0] slv0_awlen ;
wire  [2:0] slv0_awsize ;
wire  [EXTRAS-1:0] slv0_awextras ;
wire  [1:0] slv0_awburst ;
wire  slv0_awvalid ;
reg  slv0_awready ;
wire  [DWID-1:0] slv0_wdata ;
wire  [WSTRB-1:0] slv0_wstrb ;
wire  slv0_wlast ;
wire  slv0_wvalid ;
reg  slv0_wready ;
reg  [IDWID-1:0] slv0_bid ;
reg  [1:0] slv0_bresp ;
reg  slv0_bvalid ;
wire  slv0_bready ;

initial slv0_arready = 0;
initial slv0_awready = 0;
initial slv0_rvalid = 0;
initial slv0_bvalid = 0;

// reg  [2:0] slv1_awsize ; initial slv1_awsize = 0;
// reg  [2:0] slv1_arsize ; initial slv1_arsize = 0;

wire  [IDWID-1:0] slv1_arid ;
wire  [31:0] slv1_araddr ;
wire  [7:0] slv1_arlen ;
wire  [2:0] slv1_arsize ;
wire  [EXTRAS-1:0] slv1_arextras ;
wire  [1:0] slv1_arburst ;
wire  slv1_arvalid ;
reg  slv1_arready ;
reg  [IDWID-1:0] slv1_rid ;
reg  [DWID-1:0] slv1_rdata ;
reg  [1:0] slv1_rresp ;
reg  slv1_rlast ;
reg  slv1_rvalid ;
wire  slv1_rready ;

wire  [IDWID-1:0] slv1_awid ;
wire  [31:0] slv1_awaddr ;
wire  [7:0] slv1_awlen ;
wire  [2:0] slv1_awsize ;
wire  [EXTRAS-1:0] slv1_awextras ;
wire  [1:0] slv1_awburst ;
wire  slv1_awvalid ;
reg  slv1_awready ;
wire  [DWID-1:0] slv1_wdata ;
wire  [WSTRB-1:0] slv1_wstrb ;
wire  slv1_wlast ;
wire  slv1_wvalid ;
reg  slv1_wready ;
reg  [IDWID-1:0] slv1_bid ;
reg  [1:0] slv1_bresp ;
reg  slv1_bvalid ;
wire  slv1_bready ;

initial slv1_arready = 0;
initial slv1_awready = 0;
initial slv1_rvalid = 0;
initial slv1_bvalid = 0;

// reg  [2:0] slv2_awsize ; initial slv2_awsize = 0;
// reg  [2:0] slv2_arsize ; initial slv2_arsize = 0;

wire  [IDWID-1:0] slv2_arid ;
wire  [31:0] slv2_araddr ;
wire  [7:0] slv2_arlen ;
wire  [2:0] slv2_arsize ;
wire  [EXTRAS-1:0] slv2_arextras ;
wire  [1:0] slv2_arburst ;
wire  slv2_arvalid ;
reg  slv2_arready ;
reg  [IDWID-1:0] slv2_rid ;
reg  [DWID-1:0] slv2_rdata ;
reg  [1:0] slv2_rresp ;
reg  slv2_rlast ;
reg  slv2_rvalid ;
wire  slv2_rready ;

wire  [IDWID-1:0] slv2_awid ;
wire  [31:0] slv2_awaddr ;
wire  [7:0] slv2_awlen ;
wire  [2:0] slv2_awsize ;
wire  [EXTRAS-1:0] slv2_awextras ;
wire  [1:0] slv2_awburst ;
wire  slv2_awvalid ;
reg  slv2_awready ;
wire  [DWID-1:0] slv2_wdata ;
wire  [WSTRB-1:0] slv2_wstrb ;
wire  slv2_wlast ;
wire  slv2_wvalid ;
reg  slv2_wready ;
reg  [IDWID-1:0] slv2_bid ;
reg  [1:0] slv2_bresp ;
reg  slv2_bvalid ;
wire  slv2_bready ;

initial slv2_arready = 0;
initial slv2_awready = 0;
initial slv2_rvalid = 0;
initial slv2_bvalid = 0;

// reg  [2:0] slv3_awsize ; initial slv3_awsize = 0;
// reg  [2:0] slv3_arsize ; initial slv3_arsize = 0;

wire  [IDWID-1:0] slv3_arid ;
wire  [31:0] slv3_araddr ;
wire  [7:0] slv3_arlen ;
wire  [2:0] slv3_arsize ;
wire  [EXTRAS-1:0] slv3_arextras ;
wire  [1:0] slv3_arburst ;
wire  slv3_arvalid ;
reg  slv3_arready ;
reg  [IDWID-1:0] slv3_rid ;
reg  [DWID-1:0] slv3_rdata ;
reg  [1:0] slv3_rresp ;
reg  slv3_rlast ;
reg  slv3_rvalid ;
wire  slv3_rready ;

wire  [IDWID-1:0] slv3_awid ;
wire  [31:0] slv3_awaddr ;
wire  [7:0] slv3_awlen ;
wire  [2:0] slv3_awsize ;
wire  [EXTRAS-1:0] slv3_awextras ;
wire  [1:0] slv3_awburst ;
wire  slv3_awvalid ;
reg  slv3_awready ;
wire  [DWID-1:0] slv3_wdata ;
wire  [WSTRB-1:0] slv3_wstrb ;
wire  slv3_wlast ;
wire  slv3_wvalid ;
reg  slv3_wready ;
reg  [IDWID-1:0] slv3_bid ;
reg  [1:0] slv3_bresp ;
reg  slv3_bvalid ;
wire  slv3_bready ;

initial slv3_arready = 0;
initial slv3_awready = 0;
initial slv3_rvalid = 0;
initial slv3_bvalid = 0;

// reg  [2:0] mst0_awsize ; initial mst0_awsize = 0;
// reg  [2:0] mst0_arsize ; initial mst0_arsize = 0;

reg  [IDWID-1:0] mst0_arid ;
reg  [31:0] mst0_araddr ;
reg  [7:0] mst0_arlen ;
reg  [2:0] mst0_arsize ;
reg  [EXTRAS-1:0] mst0_arextras ;
reg  [1:0] mst0_arburst ;
reg  mst0_arvalid ;
wire  mst0_arready ;
wire  [IDWID-1:0] mst0_rid ;
wire  [DWID-1:0] mst0_rdata ;
wire  [1:0] mst0_rresp ;
wire  mst0_rlast ;
wire  mst0_rvalid ;
reg  mst0_rready ;

reg  [IDWID-1:0] mst0_awid ;
reg  [31:0] mst0_awaddr ;
reg  [7:0] mst0_awlen ;
reg  [2:0] mst0_awsize ;
reg  [EXTRAS-1:0] mst0_awextras ;
reg  [1:0] mst0_awburst ;
reg  mst0_awvalid ;
wire  mst0_awready ;
reg  [DWID-1:0] mst0_wdata ;
reg  [WSTRB-1:0] mst0_wstrb ;
reg  mst0_wlast ;
reg  mst0_wvalid ;
wire  mst0_wready ;
wire  [IDWID-1:0] mst0_bid ;
wire  [1:0] mst0_bresp ;
wire  mst0_bvalid ;
reg  mst0_bready ;

initial mst0_bready = 0;
initial mst0_wvalid = 0;
initial mst0_arvalid = 0;
initial mst0_awvalid = 0;
initial mst0_rready = 0;

// reg  [2:0] mst1_awsize ; initial mst1_awsize = 0;
// reg  [2:0] mst1_arsize ; initial mst1_arsize = 0;

reg  [IDWID-1:0] mst1_arid ;
reg  [31:0] mst1_araddr ;
reg  [7:0] mst1_arlen ;
reg  [2:0] mst1_arsize ;
reg  [EXTRAS-1:0] mst1_arextras ;
reg  [1:0] mst1_arburst ;
reg  mst1_arvalid ;
wire  mst1_arready ;
wire  [IDWID-1:0] mst1_rid ;
wire  [DWID-1:0] mst1_rdata ;
wire  [1:0] mst1_rresp ;
wire  mst1_rlast ;
wire  mst1_rvalid ;
reg  mst1_rready ;

reg  [IDWID-1:0] mst1_awid ;
reg  [31:0] mst1_awaddr ;
reg  [7:0] mst1_awlen ;
reg  [2:0] mst1_awsize ;
reg  [EXTRAS-1:0] mst1_awextras ;
reg  [1:0] mst1_awburst ;
reg  mst1_awvalid ;
wire  mst1_awready ;
reg  [DWID-1:0] mst1_wdata ;
reg  [WSTRB-1:0] mst1_wstrb ;
reg  mst1_wlast ;
reg  mst1_wvalid ;
wire  mst1_wready ;
wire  [IDWID-1:0] mst1_bid ;
wire  [1:0] mst1_bresp ;
wire  mst1_bvalid ;
reg  mst1_bready ;

initial mst1_bready = 0;
initial mst1_wvalid = 0;
initial mst1_arvalid = 0;
initial mst1_awvalid = 0;
initial mst1_rready = 0;

// reg  [2:0] mst10_awsize ; initial mst10_awsize = 0;
// reg  [2:0] mst10_arsize ; initial mst10_arsize = 0;

reg  [IDWID-1:0] mst10_arid ;
reg  [31:0] mst10_araddr ;
reg  [7:0] mst10_arlen ;
reg  [2:0] mst10_arsize ;
reg  [EXTRAS-1:0] mst10_arextras ;
reg  [1:0] mst10_arburst ;
reg  mst10_arvalid ;
wire  mst10_arready ;
wire  [IDWID-1:0] mst10_rid ;
wire  [DWID-1:0] mst10_rdata ;
wire  [1:0] mst10_rresp ;
wire  mst10_rlast ;
wire  mst10_rvalid ;
reg  mst10_rready ;

reg  [IDWID-1:0] mst10_awid ;
reg  [31:0] mst10_awaddr ;
reg  [7:0] mst10_awlen ;
reg  [2:0] mst10_awsize ;
reg  [EXTRAS-1:0] mst10_awextras ;
reg  [1:0] mst10_awburst ;
reg  mst10_awvalid ;
wire  mst10_awready ;
reg  [DWID-1:0] mst10_wdata ;
reg  [WSTRB-1:0] mst10_wstrb ;
reg  mst10_wlast ;
reg  mst10_wvalid ;
wire  mst10_wready ;
wire  [IDWID-1:0] mst10_bid ;
wire  [1:0] mst10_bresp ;
wire  mst10_bvalid ;
reg  mst10_bready ;

initial mst10_bready = 0;
initial mst10_wvalid = 0;
initial mst10_arvalid = 0;
initial mst10_awvalid = 0;
initial mst10_rready = 0;

// reg  [2:0] mst11_awsize ; initial mst11_awsize = 0;
// reg  [2:0] mst11_arsize ; initial mst11_arsize = 0;

reg  [IDWID-1:0] mst11_arid ;
reg  [31:0] mst11_araddr ;
reg  [7:0] mst11_arlen ;
reg  [2:0] mst11_arsize ;
reg  [EXTRAS-1:0] mst11_arextras ;
reg  [1:0] mst11_arburst ;
reg  mst11_arvalid ;
wire  mst11_arready ;
wire  [IDWID-1:0] mst11_rid ;
wire  [DWID-1:0] mst11_rdata ;
wire  [1:0] mst11_rresp ;
wire  mst11_rlast ;
wire  mst11_rvalid ;
reg  mst11_rready ;

reg  [IDWID-1:0] mst11_awid ;
reg  [31:0] mst11_awaddr ;
reg  [7:0] mst11_awlen ;
reg  [2:0] mst11_awsize ;
reg  [EXTRAS-1:0] mst11_awextras ;
reg  [1:0] mst11_awburst ;
reg  mst11_awvalid ;
wire  mst11_awready ;
reg  [DWID-1:0] mst11_wdata ;
reg  [WSTRB-1:0] mst11_wstrb ;
reg  mst11_wlast ;
reg  mst11_wvalid ;
wire  mst11_wready ;
wire  [IDWID-1:0] mst11_bid ;
wire  [1:0] mst11_bresp ;
wire  mst11_bvalid ;
reg  mst11_bready ;

initial mst11_bready = 0;
initial mst11_wvalid = 0;
initial mst11_arvalid = 0;
initial mst11_awvalid = 0;
initial mst11_rready = 0;

// reg  [2:0] mst12_awsize ; initial mst12_awsize = 0;
// reg  [2:0] mst12_arsize ; initial mst12_arsize = 0;

reg  [IDWID-1:0] mst12_arid ;
reg  [31:0] mst12_araddr ;
reg  [7:0] mst12_arlen ;
reg  [2:0] mst12_arsize ;
reg  [EXTRAS-1:0] mst12_arextras ;
reg  [1:0] mst12_arburst ;
reg  mst12_arvalid ;
wire  mst12_arready ;
wire  [IDWID-1:0] mst12_rid ;
wire  [DWID-1:0] mst12_rdata ;
wire  [1:0] mst12_rresp ;
wire  mst12_rlast ;
wire  mst12_rvalid ;
reg  mst12_rready ;

reg  [IDWID-1:0] mst12_awid ;
reg  [31:0] mst12_awaddr ;
reg  [7:0] mst12_awlen ;
reg  [2:0] mst12_awsize ;
reg  [EXTRAS-1:0] mst12_awextras ;
reg  [1:0] mst12_awburst ;
reg  mst12_awvalid ;
wire  mst12_awready ;
reg  [DWID-1:0] mst12_wdata ;
reg  [WSTRB-1:0] mst12_wstrb ;
reg  mst12_wlast ;
reg  mst12_wvalid ;
wire  mst12_wready ;
wire  [IDWID-1:0] mst12_bid ;
wire  [1:0] mst12_bresp ;
wire  mst12_bvalid ;
reg  mst12_bready ;

initial mst12_bready = 0;
initial mst12_wvalid = 0;
initial mst12_arvalid = 0;
initial mst12_awvalid = 0;
initial mst12_rready = 0;

// reg  [2:0] mst13_awsize ; initial mst13_awsize = 0;
// reg  [2:0] mst13_arsize ; initial mst13_arsize = 0;

reg  [IDWID-1:0] mst13_arid ;
reg  [31:0] mst13_araddr ;
reg  [7:0] mst13_arlen ;
reg  [2:0] mst13_arsize ;
reg  [EXTRAS-1:0] mst13_arextras ;
reg  [1:0] mst13_arburst ;
reg  mst13_arvalid ;
wire  mst13_arready ;
wire  [IDWID-1:0] mst13_rid ;
wire  [DWID-1:0] mst13_rdata ;
wire  [1:0] mst13_rresp ;
wire  mst13_rlast ;
wire  mst13_rvalid ;
reg  mst13_rready ;

reg  [IDWID-1:0] mst13_awid ;
reg  [31:0] mst13_awaddr ;
reg  [7:0] mst13_awlen ;
reg  [2:0] mst13_awsize ;
reg  [EXTRAS-1:0] mst13_awextras ;
reg  [1:0] mst13_awburst ;
reg  mst13_awvalid ;
wire  mst13_awready ;
reg  [DWID-1:0] mst13_wdata ;
reg  [WSTRB-1:0] mst13_wstrb ;
reg  mst13_wlast ;
reg  mst13_wvalid ;
wire  mst13_wready ;
wire  [IDWID-1:0] mst13_bid ;
wire  [1:0] mst13_bresp ;
wire  mst13_bvalid ;
reg  mst13_bready ;

initial mst13_bready = 0;
initial mst13_wvalid = 0;
initial mst13_arvalid = 0;
initial mst13_awvalid = 0;
initial mst13_rready = 0;

// reg  [2:0] mst14_awsize ; initial mst14_awsize = 0;
// reg  [2:0] mst14_arsize ; initial mst14_arsize = 0;

reg  [IDWID-1:0] mst14_arid ;
reg  [31:0] mst14_araddr ;
reg  [7:0] mst14_arlen ;
reg  [2:0] mst14_arsize ;
reg  [EXTRAS-1:0] mst14_arextras ;
reg  [1:0] mst14_arburst ;
reg  mst14_arvalid ;
wire  mst14_arready ;
wire  [IDWID-1:0] mst14_rid ;
wire  [DWID-1:0] mst14_rdata ;
wire  [1:0] mst14_rresp ;
wire  mst14_rlast ;
wire  mst14_rvalid ;
reg  mst14_rready ;

reg  [IDWID-1:0] mst14_awid ;
reg  [31:0] mst14_awaddr ;
reg  [7:0] mst14_awlen ;
reg  [2:0] mst14_awsize ;
reg  [EXTRAS-1:0] mst14_awextras ;
reg  [1:0] mst14_awburst ;
reg  mst14_awvalid ;
wire  mst14_awready ;
reg  [DWID-1:0] mst14_wdata ;
reg  [WSTRB-1:0] mst14_wstrb ;
reg  mst14_wlast ;
reg  mst14_wvalid ;
wire  mst14_wready ;
wire  [IDWID-1:0] mst14_bid ;
wire  [1:0] mst14_bresp ;
wire  mst14_bvalid ;
reg  mst14_bready ;

initial mst14_bready = 0;
initial mst14_wvalid = 0;
initial mst14_arvalid = 0;
initial mst14_awvalid = 0;
initial mst14_rready = 0;

// reg  [2:0] mst15_awsize ; initial mst15_awsize = 0;
// reg  [2:0] mst15_arsize ; initial mst15_arsize = 0;

reg  [IDWID-1:0] mst15_arid ;
reg  [31:0] mst15_araddr ;
reg  [7:0] mst15_arlen ;
reg  [2:0] mst15_arsize ;
reg  [EXTRAS-1:0] mst15_arextras ;
reg  [1:0] mst15_arburst ;
reg  mst15_arvalid ;
wire  mst15_arready ;
wire  [IDWID-1:0] mst15_rid ;
wire  [DWID-1:0] mst15_rdata ;
wire  [1:0] mst15_rresp ;
wire  mst15_rlast ;
wire  mst15_rvalid ;
reg  mst15_rready ;

reg  [IDWID-1:0] mst15_awid ;
reg  [31:0] mst15_awaddr ;
reg  [7:0] mst15_awlen ;
reg  [2:0] mst15_awsize ;
reg  [EXTRAS-1:0] mst15_awextras ;
reg  [1:0] mst15_awburst ;
reg  mst15_awvalid ;
wire  mst15_awready ;
reg  [DWID-1:0] mst15_wdata ;
reg  [WSTRB-1:0] mst15_wstrb ;
reg  mst15_wlast ;
reg  mst15_wvalid ;
wire  mst15_wready ;
wire  [IDWID-1:0] mst15_bid ;
wire  [1:0] mst15_bresp ;
wire  mst15_bvalid ;
reg  mst15_bready ;

initial mst15_bready = 0;
initial mst15_wvalid = 0;
initial mst15_arvalid = 0;
initial mst15_awvalid = 0;
initial mst15_rready = 0;

// reg  [2:0] mst2_awsize ; initial mst2_awsize = 0;
// reg  [2:0] mst2_arsize ; initial mst2_arsize = 0;

reg  [IDWID-1:0] mst2_arid ;
reg  [31:0] mst2_araddr ;
reg  [7:0] mst2_arlen ;
reg  [2:0] mst2_arsize ;
reg  [EXTRAS-1:0] mst2_arextras ;
reg  [1:0] mst2_arburst ;
reg  mst2_arvalid ;
wire  mst2_arready ;
wire  [IDWID-1:0] mst2_rid ;
wire  [DWID-1:0] mst2_rdata ;
wire  [1:0] mst2_rresp ;
wire  mst2_rlast ;
wire  mst2_rvalid ;
reg  mst2_rready ;

reg  [IDWID-1:0] mst2_awid ;
reg  [31:0] mst2_awaddr ;
reg  [7:0] mst2_awlen ;
reg  [2:0] mst2_awsize ;
reg  [EXTRAS-1:0] mst2_awextras ;
reg  [1:0] mst2_awburst ;
reg  mst2_awvalid ;
wire  mst2_awready ;
reg  [DWID-1:0] mst2_wdata ;
reg  [WSTRB-1:0] mst2_wstrb ;
reg  mst2_wlast ;
reg  mst2_wvalid ;
wire  mst2_wready ;
wire  [IDWID-1:0] mst2_bid ;
wire  [1:0] mst2_bresp ;
wire  mst2_bvalid ;
reg  mst2_bready ;

initial mst2_bready = 0;
initial mst2_wvalid = 0;
initial mst2_arvalid = 0;
initial mst2_awvalid = 0;
initial mst2_rready = 0;

// reg  [2:0] mst3_awsize ; initial mst3_awsize = 0;
// reg  [2:0] mst3_arsize ; initial mst3_arsize = 0;

reg  [IDWID-1:0] mst3_arid ;
reg  [31:0] mst3_araddr ;
reg  [7:0] mst3_arlen ;
reg  [2:0] mst3_arsize ;
reg  [EXTRAS-1:0] mst3_arextras ;
reg  [1:0] mst3_arburst ;
reg  mst3_arvalid ;
wire  mst3_arready ;
wire  [IDWID-1:0] mst3_rid ;
wire  [DWID-1:0] mst3_rdata ;
wire  [1:0] mst3_rresp ;
wire  mst3_rlast ;
wire  mst3_rvalid ;
reg  mst3_rready ;

reg  [IDWID-1:0] mst3_awid ;
reg  [31:0] mst3_awaddr ;
reg  [7:0] mst3_awlen ;
reg  [2:0] mst3_awsize ;
reg  [EXTRAS-1:0] mst3_awextras ;
reg  [1:0] mst3_awburst ;
reg  mst3_awvalid ;
wire  mst3_awready ;
reg  [DWID-1:0] mst3_wdata ;
reg  [WSTRB-1:0] mst3_wstrb ;
reg  mst3_wlast ;
reg  mst3_wvalid ;
wire  mst3_wready ;
wire  [IDWID-1:0] mst3_bid ;
wire  [1:0] mst3_bresp ;
wire  mst3_bvalid ;
reg  mst3_bready ;

initial mst3_bready = 0;
initial mst3_wvalid = 0;
initial mst3_arvalid = 0;
initial mst3_awvalid = 0;
initial mst3_rready = 0;

// reg  [2:0] mst4_awsize ; initial mst4_awsize = 0;
// reg  [2:0] mst4_arsize ; initial mst4_arsize = 0;

reg  [IDWID-1:0] mst4_arid ;
reg  [31:0] mst4_araddr ;
reg  [7:0] mst4_arlen ;
reg  [2:0] mst4_arsize ;
reg  [EXTRAS-1:0] mst4_arextras ;
reg  [1:0] mst4_arburst ;
reg  mst4_arvalid ;
wire  mst4_arready ;
wire  [IDWID-1:0] mst4_rid ;
wire  [DWID-1:0] mst4_rdata ;
wire  [1:0] mst4_rresp ;
wire  mst4_rlast ;
wire  mst4_rvalid ;
reg  mst4_rready ;

reg  [IDWID-1:0] mst4_awid ;
reg  [31:0] mst4_awaddr ;
reg  [7:0] mst4_awlen ;
reg  [2:0] mst4_awsize ;
reg  [EXTRAS-1:0] mst4_awextras ;
reg  [1:0] mst4_awburst ;
reg  mst4_awvalid ;
wire  mst4_awready ;
reg  [DWID-1:0] mst4_wdata ;
reg  [WSTRB-1:0] mst4_wstrb ;
reg  mst4_wlast ;
reg  mst4_wvalid ;
wire  mst4_wready ;
wire  [IDWID-1:0] mst4_bid ;
wire  [1:0] mst4_bresp ;
wire  mst4_bvalid ;
reg  mst4_bready ;

initial mst4_bready = 0;
initial mst4_wvalid = 0;
initial mst4_arvalid = 0;
initial mst4_awvalid = 0;
initial mst4_rready = 0;

// reg  [2:0] mst5_awsize ; initial mst5_awsize = 0;
// reg  [2:0] mst5_arsize ; initial mst5_arsize = 0;

reg  [IDWID-1:0] mst5_arid ;
reg  [31:0] mst5_araddr ;
reg  [7:0] mst5_arlen ;
reg  [2:0] mst5_arsize ;
reg  [EXTRAS-1:0] mst5_arextras ;
reg  [1:0] mst5_arburst ;
reg  mst5_arvalid ;
wire  mst5_arready ;
wire  [IDWID-1:0] mst5_rid ;
wire  [DWID-1:0] mst5_rdata ;
wire  [1:0] mst5_rresp ;
wire  mst5_rlast ;
wire  mst5_rvalid ;
reg  mst5_rready ;

reg  [IDWID-1:0] mst5_awid ;
reg  [31:0] mst5_awaddr ;
reg  [7:0] mst5_awlen ;
reg  [2:0] mst5_awsize ;
reg  [EXTRAS-1:0] mst5_awextras ;
reg  [1:0] mst5_awburst ;
reg  mst5_awvalid ;
wire  mst5_awready ;
reg  [DWID-1:0] mst5_wdata ;
reg  [WSTRB-1:0] mst5_wstrb ;
reg  mst5_wlast ;
reg  mst5_wvalid ;
wire  mst5_wready ;
wire  [IDWID-1:0] mst5_bid ;
wire  [1:0] mst5_bresp ;
wire  mst5_bvalid ;
reg  mst5_bready ;

initial mst5_bready = 0;
initial mst5_wvalid = 0;
initial mst5_arvalid = 0;
initial mst5_awvalid = 0;
initial mst5_rready = 0;

// reg  [2:0] mst6_awsize ; initial mst6_awsize = 0;
// reg  [2:0] mst6_arsize ; initial mst6_arsize = 0;

reg  [IDWID-1:0] mst6_arid ;
reg  [31:0] mst6_araddr ;
reg  [7:0] mst6_arlen ;
reg  [2:0] mst6_arsize ;
reg  [EXTRAS-1:0] mst6_arextras ;
reg  [1:0] mst6_arburst ;
reg  mst6_arvalid ;
wire  mst6_arready ;
wire  [IDWID-1:0] mst6_rid ;
wire  [DWID-1:0] mst6_rdata ;
wire  [1:0] mst6_rresp ;
wire  mst6_rlast ;
wire  mst6_rvalid ;
reg  mst6_rready ;

reg  [IDWID-1:0] mst6_awid ;
reg  [31:0] mst6_awaddr ;
reg  [7:0] mst6_awlen ;
reg  [2:0] mst6_awsize ;
reg  [EXTRAS-1:0] mst6_awextras ;
reg  [1:0] mst6_awburst ;
reg  mst6_awvalid ;
wire  mst6_awready ;
reg  [DWID-1:0] mst6_wdata ;
reg  [WSTRB-1:0] mst6_wstrb ;
reg  mst6_wlast ;
reg  mst6_wvalid ;
wire  mst6_wready ;
wire  [IDWID-1:0] mst6_bid ;
wire  [1:0] mst6_bresp ;
wire  mst6_bvalid ;
reg  mst6_bready ;

initial mst6_bready = 0;
initial mst6_wvalid = 0;
initial mst6_arvalid = 0;
initial mst6_awvalid = 0;
initial mst6_rready = 0;

// reg  [2:0] mst7_awsize ; initial mst7_awsize = 0;
// reg  [2:0] mst7_arsize ; initial mst7_arsize = 0;

reg  [IDWID-1:0] mst7_arid ;
reg  [31:0] mst7_araddr ;
reg  [7:0] mst7_arlen ;
reg  [2:0] mst7_arsize ;
reg  [EXTRAS-1:0] mst7_arextras ;
reg  [1:0] mst7_arburst ;
reg  mst7_arvalid ;
wire  mst7_arready ;
wire  [IDWID-1:0] mst7_rid ;
wire  [DWID-1:0] mst7_rdata ;
wire  [1:0] mst7_rresp ;
wire  mst7_rlast ;
wire  mst7_rvalid ;
reg  mst7_rready ;

reg  [IDWID-1:0] mst7_awid ;
reg  [31:0] mst7_awaddr ;
reg  [7:0] mst7_awlen ;
reg  [2:0] mst7_awsize ;
reg  [EXTRAS-1:0] mst7_awextras ;
reg  [1:0] mst7_awburst ;
reg  mst7_awvalid ;
wire  mst7_awready ;
reg  [DWID-1:0] mst7_wdata ;
reg  [WSTRB-1:0] mst7_wstrb ;
reg  mst7_wlast ;
reg  mst7_wvalid ;
wire  mst7_wready ;
wire  [IDWID-1:0] mst7_bid ;
wire  [1:0] mst7_bresp ;
wire  mst7_bvalid ;
reg  mst7_bready ;

initial mst7_bready = 0;
initial mst7_wvalid = 0;
initial mst7_arvalid = 0;
initial mst7_awvalid = 0;
initial mst7_rready = 0;

// reg  [2:0] mst8_awsize ; initial mst8_awsize = 0;
// reg  [2:0] mst8_arsize ; initial mst8_arsize = 0;

reg  [IDWID-1:0] mst8_arid ;
reg  [31:0] mst8_araddr ;
reg  [7:0] mst8_arlen ;
reg  [2:0] mst8_arsize ;
reg  [EXTRAS-1:0] mst8_arextras ;
reg  [1:0] mst8_arburst ;
reg  mst8_arvalid ;
wire  mst8_arready ;
wire  [IDWID-1:0] mst8_rid ;
wire  [DWID-1:0] mst8_rdata ;
wire  [1:0] mst8_rresp ;
wire  mst8_rlast ;
wire  mst8_rvalid ;
reg  mst8_rready ;

reg  [IDWID-1:0] mst8_awid ;
reg  [31:0] mst8_awaddr ;
reg  [7:0] mst8_awlen ;
reg  [2:0] mst8_awsize ;
reg  [EXTRAS-1:0] mst8_awextras ;
reg  [1:0] mst8_awburst ;
reg  mst8_awvalid ;
wire  mst8_awready ;
reg  [DWID-1:0] mst8_wdata ;
reg  [WSTRB-1:0] mst8_wstrb ;
reg  mst8_wlast ;
reg  mst8_wvalid ;
wire  mst8_wready ;
wire  [IDWID-1:0] mst8_bid ;
wire  [1:0] mst8_bresp ;
wire  mst8_bvalid ;
reg  mst8_bready ;

initial mst8_bready = 0;
initial mst8_wvalid = 0;
initial mst8_arvalid = 0;
initial mst8_awvalid = 0;
initial mst8_rready = 0;

// reg  [2:0] mst9_awsize ; initial mst9_awsize = 0;
// reg  [2:0] mst9_arsize ; initial mst9_arsize = 0;

reg  [IDWID-1:0] mst9_arid ;
reg  [31:0] mst9_araddr ;
reg  [7:0] mst9_arlen ;
reg  [2:0] mst9_arsize ;
reg  [EXTRAS-1:0] mst9_arextras ;
reg  [1:0] mst9_arburst ;
reg  mst9_arvalid ;
wire  mst9_arready ;
wire  [IDWID-1:0] mst9_rid ;
wire  [DWID-1:0] mst9_rdata ;
wire  [1:0] mst9_rresp ;
wire  mst9_rlast ;
wire  mst9_rvalid ;
reg  mst9_rready ;

reg  [IDWID-1:0] mst9_awid ;
reg  [31:0] mst9_awaddr ;
reg  [7:0] mst9_awlen ;
reg  [2:0] mst9_awsize ;
reg  [EXTRAS-1:0] mst9_awextras ;
reg  [1:0] mst9_awburst ;
reg  mst9_awvalid ;
wire  mst9_awready ;
reg  [DWID-1:0] mst9_wdata ;
reg  [WSTRB-1:0] mst9_wstrb ;
reg  mst9_wlast ;
reg  mst9_wvalid ;
wire  mst9_wready ;
wire  [IDWID-1:0] mst9_bid ;
wire  [1:0] mst9_bresp ;
wire  mst9_bvalid ;
reg  mst9_bready ;

initial mst9_bready = 0;
initial mst9_wvalid = 0;
initial mst9_arvalid = 0;
initial mst9_awvalid = 0;
initial mst9_rready = 0;
x16x4 dut ( .clk(clk),.rst_n(rst_n)

    ,.slv0_araddr(slv0_araddr[31:0])
    ,.slv0_arburst(slv0_arburst[1:0])
    ,.slv0_arextras(slv0_arextras[(EXTRAS - 1):0])
    ,.slv0_arid(slv0_arid)
    ,.slv0_arlen(slv0_arlen)
    ,.slv0_arsize(slv0_arsize)
    ,.slv0_arready(slv0_arready)
    ,.slv0_arvalid(slv0_arvalid)
    ,.slv0_awaddr(slv0_awaddr[31:0])
    ,.slv0_awburst(slv0_awburst[1:0])
    ,.slv0_awextras(slv0_awextras[(EXTRAS - 1):0])
    ,.slv0_awid(slv0_awid[(IDWID - 1):0])
    ,.slv0_awlen(slv0_awlen)
    ,.slv0_awsize(slv0_awsize)
    ,.slv0_awready(slv0_awready)
    ,.slv0_awvalid(slv0_awvalid)
    ,.slv0_bid(slv0_bid[(IDWID - 1):0])
    ,.slv0_bready(slv0_bready)
    ,.slv0_bresp(slv0_bresp[1:0])
    ,.slv0_bvalid(slv0_bvalid)
    ,.slv0_rdata(slv0_rdata[(DWID - 1):0])
    ,.slv0_rid(slv0_rid[(IDWID - 1):0])
    ,.slv0_rlast(slv0_rlast)
    ,.slv0_rready(slv0_rready)
    ,.slv0_rresp(slv0_rresp[1:0])
    ,.slv0_rvalid(slv0_rvalid)
    ,.slv0_wdata(slv0_wdata[(DWID - 1):0])
    ,.slv0_wlast(slv0_wlast)
    ,.slv0_wready(slv0_wready)
    ,.slv0_wstrb(slv0_wstrb[(WSTRB - 1):0])
    ,.slv0_wvalid(slv0_wvalid)


    ,.slv1_araddr(slv1_araddr[31:0])
    ,.slv1_arburst(slv1_arburst[1:0])
    ,.slv1_arextras(slv1_arextras[(EXTRAS - 1):0])
    ,.slv1_arid(slv1_arid)
    ,.slv1_arlen(slv1_arlen)
    ,.slv1_arsize(slv1_arsize)
    ,.slv1_arready(slv1_arready)
    ,.slv1_arvalid(slv1_arvalid)
    ,.slv1_awaddr(slv1_awaddr[31:0])
    ,.slv1_awburst(slv1_awburst[1:0])
    ,.slv1_awextras(slv1_awextras[(EXTRAS - 1):0])
    ,.slv1_awid(slv1_awid[(IDWID - 1):0])
    ,.slv1_awlen(slv1_awlen)
    ,.slv1_awsize(slv1_awsize)
    ,.slv1_awready(slv1_awready)
    ,.slv1_awvalid(slv1_awvalid)
    ,.slv1_bid(slv1_bid[(IDWID - 1):0])
    ,.slv1_bready(slv1_bready)
    ,.slv1_bresp(slv1_bresp[1:0])
    ,.slv1_bvalid(slv1_bvalid)
    ,.slv1_rdata(slv1_rdata[(DWID - 1):0])
    ,.slv1_rid(slv1_rid[(IDWID - 1):0])
    ,.slv1_rlast(slv1_rlast)
    ,.slv1_rready(slv1_rready)
    ,.slv1_rresp(slv1_rresp[1:0])
    ,.slv1_rvalid(slv1_rvalid)
    ,.slv1_wdata(slv1_wdata[(DWID - 1):0])
    ,.slv1_wlast(slv1_wlast)
    ,.slv1_wready(slv1_wready)
    ,.slv1_wstrb(slv1_wstrb[(WSTRB - 1):0])
    ,.slv1_wvalid(slv1_wvalid)


    ,.slv2_araddr(slv2_araddr[31:0])
    ,.slv2_arburst(slv2_arburst[1:0])
    ,.slv2_arextras(slv2_arextras[(EXTRAS - 1):0])
    ,.slv2_arid(slv2_arid)
    ,.slv2_arlen(slv2_arlen)
    ,.slv2_arsize(slv2_arsize)
    ,.slv2_arready(slv2_arready)
    ,.slv2_arvalid(slv2_arvalid)
    ,.slv2_awaddr(slv2_awaddr[31:0])
    ,.slv2_awburst(slv2_awburst[1:0])
    ,.slv2_awextras(slv2_awextras[(EXTRAS - 1):0])
    ,.slv2_awid(slv2_awid[(IDWID - 1):0])
    ,.slv2_awlen(slv2_awlen)
    ,.slv2_awsize(slv2_awsize)
    ,.slv2_awready(slv2_awready)
    ,.slv2_awvalid(slv2_awvalid)
    ,.slv2_bid(slv2_bid[(IDWID - 1):0])
    ,.slv2_bready(slv2_bready)
    ,.slv2_bresp(slv2_bresp[1:0])
    ,.slv2_bvalid(slv2_bvalid)
    ,.slv2_rdata(slv2_rdata[(DWID - 1):0])
    ,.slv2_rid(slv2_rid[(IDWID - 1):0])
    ,.slv2_rlast(slv2_rlast)
    ,.slv2_rready(slv2_rready)
    ,.slv2_rresp(slv2_rresp[1:0])
    ,.slv2_rvalid(slv2_rvalid)
    ,.slv2_wdata(slv2_wdata[(DWID - 1):0])
    ,.slv2_wlast(slv2_wlast)
    ,.slv2_wready(slv2_wready)
    ,.slv2_wstrb(slv2_wstrb[(WSTRB - 1):0])
    ,.slv2_wvalid(slv2_wvalid)


    ,.slv3_araddr(slv3_araddr[31:0])
    ,.slv3_arburst(slv3_arburst[1:0])
    ,.slv3_arextras(slv3_arextras[(EXTRAS - 1):0])
    ,.slv3_arid(slv3_arid)
    ,.slv3_arlen(slv3_arlen)
    ,.slv3_arsize(slv3_arsize)
    ,.slv3_arready(slv3_arready)
    ,.slv3_arvalid(slv3_arvalid)
    ,.slv3_awaddr(slv3_awaddr[31:0])
    ,.slv3_awburst(slv3_awburst[1:0])
    ,.slv3_awextras(slv3_awextras[(EXTRAS - 1):0])
    ,.slv3_awid(slv3_awid[(IDWID - 1):0])
    ,.slv3_awlen(slv3_awlen)
    ,.slv3_awsize(slv3_awsize)
    ,.slv3_awready(slv3_awready)
    ,.slv3_awvalid(slv3_awvalid)
    ,.slv3_bid(slv3_bid[(IDWID - 1):0])
    ,.slv3_bready(slv3_bready)
    ,.slv3_bresp(slv3_bresp[1:0])
    ,.slv3_bvalid(slv3_bvalid)
    ,.slv3_rdata(slv3_rdata[(DWID - 1):0])
    ,.slv3_rid(slv3_rid[(IDWID - 1):0])
    ,.slv3_rlast(slv3_rlast)
    ,.slv3_rready(slv3_rready)
    ,.slv3_rresp(slv3_rresp[1:0])
    ,.slv3_rvalid(slv3_rvalid)
    ,.slv3_wdata(slv3_wdata[(DWID - 1):0])
    ,.slv3_wlast(slv3_wlast)
    ,.slv3_wready(slv3_wready)
    ,.slv3_wstrb(slv3_wstrb[(WSTRB - 1):0])
    ,.slv3_wvalid(slv3_wvalid)


    ,.mst0_araddr(mst0_araddr[31:0])
    ,.mst0_arburst(mst0_arburst[1:0])
    ,.mst0_arextras(mst0_arextras[(EXTRAS - 1):0])
    ,.mst0_arid(mst0_arid)
    ,.mst0_arlen(mst0_arlen)
    ,.mst0_arsize(mst0_arsize)
    ,.mst0_arready(mst0_arready)
    ,.mst0_arvalid(mst0_arvalid)
    ,.mst0_awaddr(mst0_awaddr[31:0])
    ,.mst0_awburst(mst0_awburst[1:0])
    ,.mst0_awextras(mst0_awextras[(EXTRAS - 1):0])
    ,.mst0_awid(mst0_awid[(IDWID - 1):0])
    ,.mst0_awlen(mst0_awlen)
    ,.mst0_awsize(mst0_awsize)
    ,.mst0_awready(mst0_awready)
    ,.mst0_awvalid(mst0_awvalid)
    ,.mst0_bid(mst0_bid[(IDWID - 1):0])
    ,.mst0_bready(mst0_bready)
    ,.mst0_bresp(mst0_bresp[1:0])
    ,.mst0_bvalid(mst0_bvalid)
    ,.mst0_rdata(mst0_rdata[(DWID - 1):0])
    ,.mst0_rid(mst0_rid[(IDWID - 1):0])
    ,.mst0_rlast(mst0_rlast)
    ,.mst0_rready(mst0_rready)
    ,.mst0_rresp(mst0_rresp[1:0])
    ,.mst0_rvalid(mst0_rvalid)
    ,.mst0_wdata(mst0_wdata[(DWID - 1):0])
    ,.mst0_wlast(mst0_wlast)
    ,.mst0_wready(mst0_wready)
    ,.mst0_wstrb(mst0_wstrb[(WSTRB - 1):0])
    ,.mst0_wvalid(mst0_wvalid)

    ,.mst1_araddr(mst1_araddr[31:0])
    ,.mst1_arburst(mst1_arburst[1:0])
    ,.mst1_arextras(mst1_arextras[(EXTRAS - 1):0])
    ,.mst1_arid(mst1_arid)
    ,.mst1_arlen(mst1_arlen)
    ,.mst1_arsize(mst1_arsize)
    ,.mst1_arready(mst1_arready)
    ,.mst1_arvalid(mst1_arvalid)
    ,.mst1_awaddr(mst1_awaddr[31:0])
    ,.mst1_awburst(mst1_awburst[1:0])
    ,.mst1_awextras(mst1_awextras[(EXTRAS - 1):0])
    ,.mst1_awid(mst1_awid[(IDWID - 1):0])
    ,.mst1_awlen(mst1_awlen)
    ,.mst1_awsize(mst1_awsize)
    ,.mst1_awready(mst1_awready)
    ,.mst1_awvalid(mst1_awvalid)
    ,.mst1_bid(mst1_bid[(IDWID - 1):0])
    ,.mst1_bready(mst1_bready)
    ,.mst1_bresp(mst1_bresp[1:0])
    ,.mst1_bvalid(mst1_bvalid)
    ,.mst1_rdata(mst1_rdata[(DWID - 1):0])
    ,.mst1_rid(mst1_rid[(IDWID - 1):0])
    ,.mst1_rlast(mst1_rlast)
    ,.mst1_rready(mst1_rready)
    ,.mst1_rresp(mst1_rresp[1:0])
    ,.mst1_rvalid(mst1_rvalid)
    ,.mst1_wdata(mst1_wdata[(DWID - 1):0])
    ,.mst1_wlast(mst1_wlast)
    ,.mst1_wready(mst1_wready)
    ,.mst1_wstrb(mst1_wstrb[(WSTRB - 1):0])
    ,.mst1_wvalid(mst1_wvalid)

    ,.mst10_araddr(mst10_araddr[31:0])
    ,.mst10_arburst(mst10_arburst[1:0])
    ,.mst10_arextras(mst10_arextras[(EXTRAS - 1):0])
    ,.mst10_arid(mst10_arid)
    ,.mst10_arlen(mst10_arlen)
    ,.mst10_arsize(mst10_arsize)
    ,.mst10_arready(mst10_arready)
    ,.mst10_arvalid(mst10_arvalid)
    ,.mst10_awaddr(mst10_awaddr[31:0])
    ,.mst10_awburst(mst10_awburst[1:0])
    ,.mst10_awextras(mst10_awextras[(EXTRAS - 1):0])
    ,.mst10_awid(mst10_awid[(IDWID - 1):0])
    ,.mst10_awlen(mst10_awlen)
    ,.mst10_awsize(mst10_awsize)
    ,.mst10_awready(mst10_awready)
    ,.mst10_awvalid(mst10_awvalid)
    ,.mst10_bid(mst10_bid[(IDWID - 1):0])
    ,.mst10_bready(mst10_bready)
    ,.mst10_bresp(mst10_bresp[1:0])
    ,.mst10_bvalid(mst10_bvalid)
    ,.mst10_rdata(mst10_rdata[(DWID - 1):0])
    ,.mst10_rid(mst10_rid[(IDWID - 1):0])
    ,.mst10_rlast(mst10_rlast)
    ,.mst10_rready(mst10_rready)
    ,.mst10_rresp(mst10_rresp[1:0])
    ,.mst10_rvalid(mst10_rvalid)
    ,.mst10_wdata(mst10_wdata[(DWID - 1):0])
    ,.mst10_wlast(mst10_wlast)
    ,.mst10_wready(mst10_wready)
    ,.mst10_wstrb(mst10_wstrb[(WSTRB - 1):0])
    ,.mst10_wvalid(mst10_wvalid)

    ,.mst11_araddr(mst11_araddr[31:0])
    ,.mst11_arburst(mst11_arburst[1:0])
    ,.mst11_arextras(mst11_arextras[(EXTRAS - 1):0])
    ,.mst11_arid(mst11_arid)
    ,.mst11_arlen(mst11_arlen)
    ,.mst11_arsize(mst11_arsize)
    ,.mst11_arready(mst11_arready)
    ,.mst11_arvalid(mst11_arvalid)
    ,.mst11_awaddr(mst11_awaddr[31:0])
    ,.mst11_awburst(mst11_awburst[1:0])
    ,.mst11_awextras(mst11_awextras[(EXTRAS - 1):0])
    ,.mst11_awid(mst11_awid[(IDWID - 1):0])
    ,.mst11_awlen(mst11_awlen)
    ,.mst11_awsize(mst11_awsize)
    ,.mst11_awready(mst11_awready)
    ,.mst11_awvalid(mst11_awvalid)
    ,.mst11_bid(mst11_bid[(IDWID - 1):0])
    ,.mst11_bready(mst11_bready)
    ,.mst11_bresp(mst11_bresp[1:0])
    ,.mst11_bvalid(mst11_bvalid)
    ,.mst11_rdata(mst11_rdata[(DWID - 1):0])
    ,.mst11_rid(mst11_rid[(IDWID - 1):0])
    ,.mst11_rlast(mst11_rlast)
    ,.mst11_rready(mst11_rready)
    ,.mst11_rresp(mst11_rresp[1:0])
    ,.mst11_rvalid(mst11_rvalid)
    ,.mst11_wdata(mst11_wdata[(DWID - 1):0])
    ,.mst11_wlast(mst11_wlast)
    ,.mst11_wready(mst11_wready)
    ,.mst11_wstrb(mst11_wstrb[(WSTRB - 1):0])
    ,.mst11_wvalid(mst11_wvalid)

    ,.mst12_araddr(mst12_araddr[31:0])
    ,.mst12_arburst(mst12_arburst[1:0])
    ,.mst12_arextras(mst12_arextras[(EXTRAS - 1):0])
    ,.mst12_arid(mst12_arid)
    ,.mst12_arlen(mst12_arlen)
    ,.mst12_arsize(mst12_arsize)
    ,.mst12_arready(mst12_arready)
    ,.mst12_arvalid(mst12_arvalid)
    ,.mst12_awaddr(mst12_awaddr[31:0])
    ,.mst12_awburst(mst12_awburst[1:0])
    ,.mst12_awextras(mst12_awextras[(EXTRAS - 1):0])
    ,.mst12_awid(mst12_awid[(IDWID - 1):0])
    ,.mst12_awlen(mst12_awlen)
    ,.mst12_awsize(mst12_awsize)
    ,.mst12_awready(mst12_awready)
    ,.mst12_awvalid(mst12_awvalid)
    ,.mst12_bid(mst12_bid[(IDWID - 1):0])
    ,.mst12_bready(mst12_bready)
    ,.mst12_bresp(mst12_bresp[1:0])
    ,.mst12_bvalid(mst12_bvalid)
    ,.mst12_rdata(mst12_rdata[(DWID - 1):0])
    ,.mst12_rid(mst12_rid[(IDWID - 1):0])
    ,.mst12_rlast(mst12_rlast)
    ,.mst12_rready(mst12_rready)
    ,.mst12_rresp(mst12_rresp[1:0])
    ,.mst12_rvalid(mst12_rvalid)
    ,.mst12_wdata(mst12_wdata[(DWID - 1):0])
    ,.mst12_wlast(mst12_wlast)
    ,.mst12_wready(mst12_wready)
    ,.mst12_wstrb(mst12_wstrb[(WSTRB - 1):0])
    ,.mst12_wvalid(mst12_wvalid)

    ,.mst13_araddr(mst13_araddr[31:0])
    ,.mst13_arburst(mst13_arburst[1:0])
    ,.mst13_arextras(mst13_arextras[(EXTRAS - 1):0])
    ,.mst13_arid(mst13_arid)
    ,.mst13_arlen(mst13_arlen)
    ,.mst13_arsize(mst13_arsize)
    ,.mst13_arready(mst13_arready)
    ,.mst13_arvalid(mst13_arvalid)
    ,.mst13_awaddr(mst13_awaddr[31:0])
    ,.mst13_awburst(mst13_awburst[1:0])
    ,.mst13_awextras(mst13_awextras[(EXTRAS - 1):0])
    ,.mst13_awid(mst13_awid[(IDWID - 1):0])
    ,.mst13_awlen(mst13_awlen)
    ,.mst13_awsize(mst13_awsize)
    ,.mst13_awready(mst13_awready)
    ,.mst13_awvalid(mst13_awvalid)
    ,.mst13_bid(mst13_bid[(IDWID - 1):0])
    ,.mst13_bready(mst13_bready)
    ,.mst13_bresp(mst13_bresp[1:0])
    ,.mst13_bvalid(mst13_bvalid)
    ,.mst13_rdata(mst13_rdata[(DWID - 1):0])
    ,.mst13_rid(mst13_rid[(IDWID - 1):0])
    ,.mst13_rlast(mst13_rlast)
    ,.mst13_rready(mst13_rready)
    ,.mst13_rresp(mst13_rresp[1:0])
    ,.mst13_rvalid(mst13_rvalid)
    ,.mst13_wdata(mst13_wdata[(DWID - 1):0])
    ,.mst13_wlast(mst13_wlast)
    ,.mst13_wready(mst13_wready)
    ,.mst13_wstrb(mst13_wstrb[(WSTRB - 1):0])
    ,.mst13_wvalid(mst13_wvalid)

    ,.mst14_araddr(mst14_araddr[31:0])
    ,.mst14_arburst(mst14_arburst[1:0])
    ,.mst14_arextras(mst14_arextras[(EXTRAS - 1):0])
    ,.mst14_arid(mst14_arid)
    ,.mst14_arlen(mst14_arlen)
    ,.mst14_arsize(mst14_arsize)
    ,.mst14_arready(mst14_arready)
    ,.mst14_arvalid(mst14_arvalid)
    ,.mst14_awaddr(mst14_awaddr[31:0])
    ,.mst14_awburst(mst14_awburst[1:0])
    ,.mst14_awextras(mst14_awextras[(EXTRAS - 1):0])
    ,.mst14_awid(mst14_awid[(IDWID - 1):0])
    ,.mst14_awlen(mst14_awlen)
    ,.mst14_awsize(mst14_awsize)
    ,.mst14_awready(mst14_awready)
    ,.mst14_awvalid(mst14_awvalid)
    ,.mst14_bid(mst14_bid[(IDWID - 1):0])
    ,.mst14_bready(mst14_bready)
    ,.mst14_bresp(mst14_bresp[1:0])
    ,.mst14_bvalid(mst14_bvalid)
    ,.mst14_rdata(mst14_rdata[(DWID - 1):0])
    ,.mst14_rid(mst14_rid[(IDWID - 1):0])
    ,.mst14_rlast(mst14_rlast)
    ,.mst14_rready(mst14_rready)
    ,.mst14_rresp(mst14_rresp[1:0])
    ,.mst14_rvalid(mst14_rvalid)
    ,.mst14_wdata(mst14_wdata[(DWID - 1):0])
    ,.mst14_wlast(mst14_wlast)
    ,.mst14_wready(mst14_wready)
    ,.mst14_wstrb(mst14_wstrb[(WSTRB - 1):0])
    ,.mst14_wvalid(mst14_wvalid)

    ,.mst15_araddr(mst15_araddr[31:0])
    ,.mst15_arburst(mst15_arburst[1:0])
    ,.mst15_arextras(mst15_arextras[(EXTRAS - 1):0])
    ,.mst15_arid(mst15_arid)
    ,.mst15_arlen(mst15_arlen)
    ,.mst15_arsize(mst15_arsize)
    ,.mst15_arready(mst15_arready)
    ,.mst15_arvalid(mst15_arvalid)
    ,.mst15_awaddr(mst15_awaddr[31:0])
    ,.mst15_awburst(mst15_awburst[1:0])
    ,.mst15_awextras(mst15_awextras[(EXTRAS - 1):0])
    ,.mst15_awid(mst15_awid[(IDWID - 1):0])
    ,.mst15_awlen(mst15_awlen)
    ,.mst15_awsize(mst15_awsize)
    ,.mst15_awready(mst15_awready)
    ,.mst15_awvalid(mst15_awvalid)
    ,.mst15_bid(mst15_bid[(IDWID - 1):0])
    ,.mst15_bready(mst15_bready)
    ,.mst15_bresp(mst15_bresp[1:0])
    ,.mst15_bvalid(mst15_bvalid)
    ,.mst15_rdata(mst15_rdata[(DWID - 1):0])
    ,.mst15_rid(mst15_rid[(IDWID - 1):0])
    ,.mst15_rlast(mst15_rlast)
    ,.mst15_rready(mst15_rready)
    ,.mst15_rresp(mst15_rresp[1:0])
    ,.mst15_rvalid(mst15_rvalid)
    ,.mst15_wdata(mst15_wdata[(DWID - 1):0])
    ,.mst15_wlast(mst15_wlast)
    ,.mst15_wready(mst15_wready)
    ,.mst15_wstrb(mst15_wstrb[(WSTRB - 1):0])
    ,.mst15_wvalid(mst15_wvalid)

    ,.mst2_araddr(mst2_araddr[31:0])
    ,.mst2_arburst(mst2_arburst[1:0])
    ,.mst2_arextras(mst2_arextras[(EXTRAS - 1):0])
    ,.mst2_arid(mst2_arid)
    ,.mst2_arlen(mst2_arlen)
    ,.mst2_arsize(mst2_arsize)
    ,.mst2_arready(mst2_arready)
    ,.mst2_arvalid(mst2_arvalid)
    ,.mst2_awaddr(mst2_awaddr[31:0])
    ,.mst2_awburst(mst2_awburst[1:0])
    ,.mst2_awextras(mst2_awextras[(EXTRAS - 1):0])
    ,.mst2_awid(mst2_awid[(IDWID - 1):0])
    ,.mst2_awlen(mst2_awlen)
    ,.mst2_awsize(mst2_awsize)
    ,.mst2_awready(mst2_awready)
    ,.mst2_awvalid(mst2_awvalid)
    ,.mst2_bid(mst2_bid[(IDWID - 1):0])
    ,.mst2_bready(mst2_bready)
    ,.mst2_bresp(mst2_bresp[1:0])
    ,.mst2_bvalid(mst2_bvalid)
    ,.mst2_rdata(mst2_rdata[(DWID - 1):0])
    ,.mst2_rid(mst2_rid[(IDWID - 1):0])
    ,.mst2_rlast(mst2_rlast)
    ,.mst2_rready(mst2_rready)
    ,.mst2_rresp(mst2_rresp[1:0])
    ,.mst2_rvalid(mst2_rvalid)
    ,.mst2_wdata(mst2_wdata[(DWID - 1):0])
    ,.mst2_wlast(mst2_wlast)
    ,.mst2_wready(mst2_wready)
    ,.mst2_wstrb(mst2_wstrb[(WSTRB - 1):0])
    ,.mst2_wvalid(mst2_wvalid)

    ,.mst3_araddr(mst3_araddr[31:0])
    ,.mst3_arburst(mst3_arburst[1:0])
    ,.mst3_arextras(mst3_arextras[(EXTRAS - 1):0])
    ,.mst3_arid(mst3_arid)
    ,.mst3_arlen(mst3_arlen)
    ,.mst3_arsize(mst3_arsize)
    ,.mst3_arready(mst3_arready)
    ,.mst3_arvalid(mst3_arvalid)
    ,.mst3_awaddr(mst3_awaddr[31:0])
    ,.mst3_awburst(mst3_awburst[1:0])
    ,.mst3_awextras(mst3_awextras[(EXTRAS - 1):0])
    ,.mst3_awid(mst3_awid[(IDWID - 1):0])
    ,.mst3_awlen(mst3_awlen)
    ,.mst3_awsize(mst3_awsize)
    ,.mst3_awready(mst3_awready)
    ,.mst3_awvalid(mst3_awvalid)
    ,.mst3_bid(mst3_bid[(IDWID - 1):0])
    ,.mst3_bready(mst3_bready)
    ,.mst3_bresp(mst3_bresp[1:0])
    ,.mst3_bvalid(mst3_bvalid)
    ,.mst3_rdata(mst3_rdata[(DWID - 1):0])
    ,.mst3_rid(mst3_rid[(IDWID - 1):0])
    ,.mst3_rlast(mst3_rlast)
    ,.mst3_rready(mst3_rready)
    ,.mst3_rresp(mst3_rresp[1:0])
    ,.mst3_rvalid(mst3_rvalid)
    ,.mst3_wdata(mst3_wdata[(DWID - 1):0])
    ,.mst3_wlast(mst3_wlast)
    ,.mst3_wready(mst3_wready)
    ,.mst3_wstrb(mst3_wstrb[(WSTRB - 1):0])
    ,.mst3_wvalid(mst3_wvalid)

    ,.mst4_araddr(mst4_araddr[31:0])
    ,.mst4_arburst(mst4_arburst[1:0])
    ,.mst4_arextras(mst4_arextras[(EXTRAS - 1):0])
    ,.mst4_arid(mst4_arid)
    ,.mst4_arlen(mst4_arlen)
    ,.mst4_arsize(mst4_arsize)
    ,.mst4_arready(mst4_arready)
    ,.mst4_arvalid(mst4_arvalid)
    ,.mst4_awaddr(mst4_awaddr[31:0])
    ,.mst4_awburst(mst4_awburst[1:0])
    ,.mst4_awextras(mst4_awextras[(EXTRAS - 1):0])
    ,.mst4_awid(mst4_awid[(IDWID - 1):0])
    ,.mst4_awlen(mst4_awlen)
    ,.mst4_awsize(mst4_awsize)
    ,.mst4_awready(mst4_awready)
    ,.mst4_awvalid(mst4_awvalid)
    ,.mst4_bid(mst4_bid[(IDWID - 1):0])
    ,.mst4_bready(mst4_bready)
    ,.mst4_bresp(mst4_bresp[1:0])
    ,.mst4_bvalid(mst4_bvalid)
    ,.mst4_rdata(mst4_rdata[(DWID - 1):0])
    ,.mst4_rid(mst4_rid[(IDWID - 1):0])
    ,.mst4_rlast(mst4_rlast)
    ,.mst4_rready(mst4_rready)
    ,.mst4_rresp(mst4_rresp[1:0])
    ,.mst4_rvalid(mst4_rvalid)
    ,.mst4_wdata(mst4_wdata[(DWID - 1):0])
    ,.mst4_wlast(mst4_wlast)
    ,.mst4_wready(mst4_wready)
    ,.mst4_wstrb(mst4_wstrb[(WSTRB - 1):0])
    ,.mst4_wvalid(mst4_wvalid)

    ,.mst5_araddr(mst5_araddr[31:0])
    ,.mst5_arburst(mst5_arburst[1:0])
    ,.mst5_arextras(mst5_arextras[(EXTRAS - 1):0])
    ,.mst5_arid(mst5_arid)
    ,.mst5_arlen(mst5_arlen)
    ,.mst5_arsize(mst5_arsize)
    ,.mst5_arready(mst5_arready)
    ,.mst5_arvalid(mst5_arvalid)
    ,.mst5_awaddr(mst5_awaddr[31:0])
    ,.mst5_awburst(mst5_awburst[1:0])
    ,.mst5_awextras(mst5_awextras[(EXTRAS - 1):0])
    ,.mst5_awid(mst5_awid[(IDWID - 1):0])
    ,.mst5_awlen(mst5_awlen)
    ,.mst5_awsize(mst5_awsize)
    ,.mst5_awready(mst5_awready)
    ,.mst5_awvalid(mst5_awvalid)
    ,.mst5_bid(mst5_bid[(IDWID - 1):0])
    ,.mst5_bready(mst5_bready)
    ,.mst5_bresp(mst5_bresp[1:0])
    ,.mst5_bvalid(mst5_bvalid)
    ,.mst5_rdata(mst5_rdata[(DWID - 1):0])
    ,.mst5_rid(mst5_rid[(IDWID - 1):0])
    ,.mst5_rlast(mst5_rlast)
    ,.mst5_rready(mst5_rready)
    ,.mst5_rresp(mst5_rresp[1:0])
    ,.mst5_rvalid(mst5_rvalid)
    ,.mst5_wdata(mst5_wdata[(DWID - 1):0])
    ,.mst5_wlast(mst5_wlast)
    ,.mst5_wready(mst5_wready)
    ,.mst5_wstrb(mst5_wstrb[(WSTRB - 1):0])
    ,.mst5_wvalid(mst5_wvalid)

    ,.mst6_araddr(mst6_araddr[31:0])
    ,.mst6_arburst(mst6_arburst[1:0])
    ,.mst6_arextras(mst6_arextras[(EXTRAS - 1):0])
    ,.mst6_arid(mst6_arid)
    ,.mst6_arlen(mst6_arlen)
    ,.mst6_arsize(mst6_arsize)
    ,.mst6_arready(mst6_arready)
    ,.mst6_arvalid(mst6_arvalid)
    ,.mst6_awaddr(mst6_awaddr[31:0])
    ,.mst6_awburst(mst6_awburst[1:0])
    ,.mst6_awextras(mst6_awextras[(EXTRAS - 1):0])
    ,.mst6_awid(mst6_awid[(IDWID - 1):0])
    ,.mst6_awlen(mst6_awlen)
    ,.mst6_awsize(mst6_awsize)
    ,.mst6_awready(mst6_awready)
    ,.mst6_awvalid(mst6_awvalid)
    ,.mst6_bid(mst6_bid[(IDWID - 1):0])
    ,.mst6_bready(mst6_bready)
    ,.mst6_bresp(mst6_bresp[1:0])
    ,.mst6_bvalid(mst6_bvalid)
    ,.mst6_rdata(mst6_rdata[(DWID - 1):0])
    ,.mst6_rid(mst6_rid[(IDWID - 1):0])
    ,.mst6_rlast(mst6_rlast)
    ,.mst6_rready(mst6_rready)
    ,.mst6_rresp(mst6_rresp[1:0])
    ,.mst6_rvalid(mst6_rvalid)
    ,.mst6_wdata(mst6_wdata[(DWID - 1):0])
    ,.mst6_wlast(mst6_wlast)
    ,.mst6_wready(mst6_wready)
    ,.mst6_wstrb(mst6_wstrb[(WSTRB - 1):0])
    ,.mst6_wvalid(mst6_wvalid)

    ,.mst7_araddr(mst7_araddr[31:0])
    ,.mst7_arburst(mst7_arburst[1:0])
    ,.mst7_arextras(mst7_arextras[(EXTRAS - 1):0])
    ,.mst7_arid(mst7_arid)
    ,.mst7_arlen(mst7_arlen)
    ,.mst7_arsize(mst7_arsize)
    ,.mst7_arready(mst7_arready)
    ,.mst7_arvalid(mst7_arvalid)
    ,.mst7_awaddr(mst7_awaddr[31:0])
    ,.mst7_awburst(mst7_awburst[1:0])
    ,.mst7_awextras(mst7_awextras[(EXTRAS - 1):0])
    ,.mst7_awid(mst7_awid[(IDWID - 1):0])
    ,.mst7_awlen(mst7_awlen)
    ,.mst7_awsize(mst7_awsize)
    ,.mst7_awready(mst7_awready)
    ,.mst7_awvalid(mst7_awvalid)
    ,.mst7_bid(mst7_bid[(IDWID - 1):0])
    ,.mst7_bready(mst7_bready)
    ,.mst7_bresp(mst7_bresp[1:0])
    ,.mst7_bvalid(mst7_bvalid)
    ,.mst7_rdata(mst7_rdata[(DWID - 1):0])
    ,.mst7_rid(mst7_rid[(IDWID - 1):0])
    ,.mst7_rlast(mst7_rlast)
    ,.mst7_rready(mst7_rready)
    ,.mst7_rresp(mst7_rresp[1:0])
    ,.mst7_rvalid(mst7_rvalid)
    ,.mst7_wdata(mst7_wdata[(DWID - 1):0])
    ,.mst7_wlast(mst7_wlast)
    ,.mst7_wready(mst7_wready)
    ,.mst7_wstrb(mst7_wstrb[(WSTRB - 1):0])
    ,.mst7_wvalid(mst7_wvalid)

    ,.mst8_araddr(mst8_araddr[31:0])
    ,.mst8_arburst(mst8_arburst[1:0])
    ,.mst8_arextras(mst8_arextras[(EXTRAS - 1):0])
    ,.mst8_arid(mst8_arid)
    ,.mst8_arlen(mst8_arlen)
    ,.mst8_arsize(mst8_arsize)
    ,.mst8_arready(mst8_arready)
    ,.mst8_arvalid(mst8_arvalid)
    ,.mst8_awaddr(mst8_awaddr[31:0])
    ,.mst8_awburst(mst8_awburst[1:0])
    ,.mst8_awextras(mst8_awextras[(EXTRAS - 1):0])
    ,.mst8_awid(mst8_awid[(IDWID - 1):0])
    ,.mst8_awlen(mst8_awlen)
    ,.mst8_awsize(mst8_awsize)
    ,.mst8_awready(mst8_awready)
    ,.mst8_awvalid(mst8_awvalid)
    ,.mst8_bid(mst8_bid[(IDWID - 1):0])
    ,.mst8_bready(mst8_bready)
    ,.mst8_bresp(mst8_bresp[1:0])
    ,.mst8_bvalid(mst8_bvalid)
    ,.mst8_rdata(mst8_rdata[(DWID - 1):0])
    ,.mst8_rid(mst8_rid[(IDWID - 1):0])
    ,.mst8_rlast(mst8_rlast)
    ,.mst8_rready(mst8_rready)
    ,.mst8_rresp(mst8_rresp[1:0])
    ,.mst8_rvalid(mst8_rvalid)
    ,.mst8_wdata(mst8_wdata[(DWID - 1):0])
    ,.mst8_wlast(mst8_wlast)
    ,.mst8_wready(mst8_wready)
    ,.mst8_wstrb(mst8_wstrb[(WSTRB - 1):0])
    ,.mst8_wvalid(mst8_wvalid)

    ,.mst9_araddr(mst9_araddr[31:0])
    ,.mst9_arburst(mst9_arburst[1:0])
    ,.mst9_arextras(mst9_arextras[(EXTRAS - 1):0])
    ,.mst9_arid(mst9_arid)
    ,.mst9_arlen(mst9_arlen)
    ,.mst9_arsize(mst9_arsize)
    ,.mst9_arready(mst9_arready)
    ,.mst9_arvalid(mst9_arvalid)
    ,.mst9_awaddr(mst9_awaddr[31:0])
    ,.mst9_awburst(mst9_awburst[1:0])
    ,.mst9_awextras(mst9_awextras[(EXTRAS - 1):0])
    ,.mst9_awid(mst9_awid[(IDWID - 1):0])
    ,.mst9_awlen(mst9_awlen)
    ,.mst9_awsize(mst9_awsize)
    ,.mst9_awready(mst9_awready)
    ,.mst9_awvalid(mst9_awvalid)
    ,.mst9_bid(mst9_bid[(IDWID - 1):0])
    ,.mst9_bready(mst9_bready)
    ,.mst9_bresp(mst9_bresp[1:0])
    ,.mst9_bvalid(mst9_bvalid)
    ,.mst9_rdata(mst9_rdata[(DWID - 1):0])
    ,.mst9_rid(mst9_rid[(IDWID - 1):0])
    ,.mst9_rlast(mst9_rlast)
    ,.mst9_rready(mst9_rready)
    ,.mst9_rresp(mst9_rresp[1:0])
    ,.mst9_rvalid(mst9_rvalid)
    ,.mst9_wdata(mst9_wdata[(DWID - 1):0])
    ,.mst9_wlast(mst9_wlast)
    ,.mst9_wready(mst9_wready)
    ,.mst9_wstrb(mst9_wstrb[(WSTRB - 1):0])
    ,.mst9_wvalid(mst9_wvalid)
);


reg [1023:0] testname;
initial begin
   if ($value$plusargs("LOG=%s",testname)) begin 
        $python("pymonname()",testname);
    end  


    if ($value$plusargs("SEQ=%s",testname)) begin 
         $display(" Running SEQ= %s.",testname); 
    end else begin
        testname = 0; 
        $display(" default test");
    end  
    #10; 
    if (testname!=0) $python("sequence()",testname);
end 
endmodule

