module atan_table_till_32k(input [9:0] addr,output [24:0] result,output [24:0] lastone);
assign result = 
    (addr==0) ? 24681426 :   //   in=10.000000 val=1.471128
    (addr==1) ? 24686601 :   //   in=10.031250 val=1.471436
    (addr==2) ? 24691744 :   //   in=10.062500 val=1.471743
    (addr==3) ? 24696856 :   //   in=10.093750 val=1.472047
    (addr==4) ? 24701936 :   //   in=10.125000 val=1.472350
    (addr==5) ? 24706986 :   //   in=10.156250 val=1.472651
    (addr==6) ? 24712004 :   //   in=10.187500 val=1.472950
    (addr==7) ? 24716993 :   //   in=10.218750 val=1.473248
    (addr==8) ? 24721951 :   //   in=10.250000 val=1.473543
    (addr==9) ? 24726879 :   //   in=10.281250 val=1.473837
    (addr==10) ? 24731778 :   //   in=10.312500 val=1.474129
    (addr==11) ? 24736647 :   //   in=10.343750 val=1.474419
    (addr==12) ? 24741488 :   //   in=10.375000 val=1.474708
    (addr==13) ? 24746299 :   //   in=10.406250 val=1.474994
    (addr==14) ? 24751082 :   //   in=10.437500 val=1.475279
    (addr==15) ? 24755837 :   //   in=10.468750 val=1.475563
    (addr==16) ? 24760563 :   //   in=10.500000 val=1.475845
    (addr==17) ? 24765262 :   //   in=10.531250 val=1.476125
    (addr==18) ? 24769934 :   //   in=10.562500 val=1.476403
    (addr==19) ? 24774578 :   //   in=10.593750 val=1.476680
    (addr==20) ? 24779194 :   //   in=10.625000 val=1.476955
    (addr==21) ? 24783785 :   //   in=10.656250 val=1.477229
    (addr==22) ? 24788348 :   //   in=10.687500 val=1.477501
    (addr==23) ? 24792885 :   //   in=10.718750 val=1.477771
    (addr==24) ? 24797396 :   //   in=10.750000 val=1.478040
    (addr==25) ? 24801881 :   //   in=10.781250 val=1.478307
    (addr==26) ? 24806340 :   //   in=10.812500 val=1.478573
    (addr==27) ? 24810774 :   //   in=10.843750 val=1.478837
    (addr==28) ? 24815183 :   //   in=10.875000 val=1.479100
    (addr==29) ? 24819566 :   //   in=10.906250 val=1.479361
    (addr==30) ? 24823925 :   //   in=10.937500 val=1.479621
    (addr==31) ? 24828259 :   //   in=10.968750 val=1.479880
    (addr==32) ? 24832568 :   //   in=11.000000 val=1.480136
    (addr==33) ? 24836854 :   //   in=11.031250 val=1.480392
    (addr==34) ? 24841115 :   //   in=11.062500 val=1.480646
    (addr==35) ? 24845353 :   //   in=11.093750 val=1.480898
    (addr==36) ? 24849566 :   //   in=11.125000 val=1.481150
    (addr==37) ? 24853757 :   //   in=11.156250 val=1.481399
    (addr==38) ? 24857924 :   //   in=11.187500 val=1.481648
    (addr==39) ? 24862068 :   //   in=11.218750 val=1.481895
    (addr==40) ? 24866190 :   //   in=11.250000 val=1.482140
    (addr==41) ? 24870289 :   //   in=11.281250 val=1.482385
    (addr==42) ? 24874365 :   //   in=11.312500 val=1.482628
    (addr==43) ? 24878419 :   //   in=11.343750 val=1.482869
    (addr==44) ? 24882451 :   //   in=11.375000 val=1.483110
    (addr==45) ? 24886461 :   //   in=11.406250 val=1.483349
    (addr==46) ? 24890449 :   //   in=11.437500 val=1.483586
    (addr==47) ? 24894416 :   //   in=11.468750 val=1.483823
    (addr==48) ? 24898361 :   //   in=11.500000 val=1.484058
    (addr==49) ? 24902285 :   //   in=11.531250 val=1.484292
    (addr==50) ? 24906188 :   //   in=11.562500 val=1.484525
    (addr==51) ? 24910070 :   //   in=11.593750 val=1.484756
    (addr==52) ? 24913931 :   //   in=11.625000 val=1.484986
    (addr==53) ? 24917772 :   //   in=11.656250 val=1.485215
    (addr==54) ? 24921593 :   //   in=11.687500 val=1.485443
    (addr==55) ? 24925393 :   //   in=11.718750 val=1.485669
    (addr==56) ? 24929173 :   //   in=11.750000 val=1.485895
    (addr==57) ? 24932933 :   //   in=11.781250 val=1.486119
    (addr==58) ? 24936674 :   //   in=11.812500 val=1.486342
    (addr==59) ? 24940395 :   //   in=11.843750 val=1.486563
    (addr==60) ? 24944096 :   //   in=11.875000 val=1.486784
    (addr==61) ? 24947778 :   //   in=11.906250 val=1.487003
    (addr==62) ? 24951441 :   //   in=11.937500 val=1.487222
    (addr==63) ? 24955085 :   //   in=11.968750 val=1.487439
    (addr==64) ? 24958710 :   //   in=12.000000 val=1.487655
    (addr==65) ? 24962317 :   //   in=12.031250 val=1.487870
    (addr==66) ? 24965905 :   //   in=12.062500 val=1.488084
    (addr==67) ? 24969474 :   //   in=12.093750 val=1.488297
    (addr==68) ? 24973025 :   //   in=12.125000 val=1.488508
    (addr==69) ? 24976558 :   //   in=12.156250 val=1.488719
    (addr==70) ? 24980074 :   //   in=12.187500 val=1.488928
    (addr==71) ? 24983571 :   //   in=12.218750 val=1.489137
    (addr==72) ? 24987050 :   //   in=12.250000 val=1.489344
    (addr==73) ? 24990512 :   //   in=12.281250 val=1.489551
    (addr==74) ? 24993957 :   //   in=12.312500 val=1.489756
    (addr==75) ? 24997384 :   //   in=12.343750 val=1.489960
    (addr==76) ? 25000794 :   //   in=12.375000 val=1.490163
    (addr==77) ? 25004186 :   //   in=12.406250 val=1.490366
    (addr==78) ? 25007562 :   //   in=12.437500 val=1.490567
    (addr==79) ? 25010921 :   //   in=12.468750 val=1.490767
    (addr==80) ? 25014264 :   //   in=12.500000 val=1.490966
    (addr==81) ? 25017590 :   //   in=12.531250 val=1.491165
    (addr==82) ? 25020899 :   //   in=12.562500 val=1.491362
    (addr==83) ? 25024192 :   //   in=12.593750 val=1.491558
    (addr==84) ? 25027469 :   //   in=12.625000 val=1.491753
    (addr==85) ? 25030730 :   //   in=12.656250 val=1.491948
    (addr==86) ? 25033975 :   //   in=12.687500 val=1.492141
    (addr==87) ? 25037204 :   //   in=12.718750 val=1.492334
    (addr==88) ? 25040417 :   //   in=12.750000 val=1.492525
    (addr==89) ? 25043615 :   //   in=12.781250 val=1.492716
    (addr==90) ? 25046797 :   //   in=12.812500 val=1.492905
    (addr==91) ? 25049963 :   //   in=12.843750 val=1.493094
    (addr==92) ? 25053115 :   //   in=12.875000 val=1.493282
    (addr==93) ? 25056251 :   //   in=12.906250 val=1.493469
    (addr==94) ? 25059372 :   //   in=12.937500 val=1.493655
    (addr==95) ? 25062479 :   //   in=12.968750 val=1.493840
    (addr==96) ? 25065570 :   //   in=13.000000 val=1.494024
    (addr==97) ? 25068647 :   //   in=13.031250 val=1.494208
    (addr==98) ? 25071709 :   //   in=13.062500 val=1.494390
    (addr==99) ? 25074756 :   //   in=13.093750 val=1.494572
    (addr==100) ? 25077790 :   //   in=13.125000 val=1.494753
    (addr==101) ? 25080808 :   //   in=13.156250 val=1.494933
    (addr==102) ? 25083813 :   //   in=13.187500 val=1.495112
    (addr==103) ? 25086803 :   //   in=13.218750 val=1.495290
    (addr==104) ? 25089780 :   //   in=13.250000 val=1.495467
    (addr==105) ? 25092742 :   //   in=13.281250 val=1.495644
    (addr==106) ? 25095691 :   //   in=13.312500 val=1.495820
    (addr==107) ? 25098626 :   //   in=13.343750 val=1.495995
    (addr==108) ? 25101547 :   //   in=13.375000 val=1.496169
    (addr==109) ? 25104455 :   //   in=13.406250 val=1.496342
    (addr==110) ? 25107349 :   //   in=13.437500 val=1.496515
    (addr==111) ? 25110230 :   //   in=13.468750 val=1.496686
    (addr==112) ? 25113098 :   //   in=13.500000 val=1.496857
    (addr==113) ? 25115952 :   //   in=13.531250 val=1.497027
    (addr==114) ? 25118793 :   //   in=13.562500 val=1.497197
    (addr==115) ? 25121622 :   //   in=13.593750 val=1.497365
    (addr==116) ? 25124437 :   //   in=13.625000 val=1.497533
    (addr==117) ? 25127240 :   //   in=13.656250 val=1.497700
    (addr==118) ? 25130030 :   //   in=13.687500 val=1.497867
    (addr==119) ? 25132807 :   //   in=13.718750 val=1.498032
    (addr==120) ? 25135572 :   //   in=13.750000 val=1.498197
    (addr==121) ? 25138324 :   //   in=13.781250 val=1.498361
    (addr==122) ? 25141064 :   //   in=13.812500 val=1.498524
    (addr==123) ? 25143792 :   //   in=13.843750 val=1.498687
    (addr==124) ? 25146507 :   //   in=13.875000 val=1.498849
    (addr==125) ? 25149210 :   //   in=13.906250 val=1.499010
    (addr==126) ? 25151902 :   //   in=13.937500 val=1.499170
    (addr==127) ? 25154581 :   //   in=13.968750 val=1.499330
    (addr==128) ? 25157248 :   //   in=14.000000 val=1.499489
    (addr==129) ? 25159903 :   //   in=14.031250 val=1.499647
    (addr==130) ? 25162547 :   //   in=14.062500 val=1.499805
    (addr==131) ? 25165179 :   //   in=14.093750 val=1.499962
    (addr==132) ? 25167800 :   //   in=14.125000 val=1.500118
    (addr==133) ? 25170409 :   //   in=14.156250 val=1.500273
    (addr==134) ? 25173006 :   //   in=14.187500 val=1.500428
    (addr==135) ? 25175592 :   //   in=14.218750 val=1.500582
    (addr==136) ? 25178167 :   //   in=14.250000 val=1.500736
    (addr==137) ? 25180731 :   //   in=14.281250 val=1.500889
    (addr==138) ? 25183283 :   //   in=14.312500 val=1.501041
    (addr==139) ? 25185825 :   //   in=14.343750 val=1.501192
    (addr==140) ? 25188355 :   //   in=14.375000 val=1.501343
    (addr==141) ? 25190875 :   //   in=14.406250 val=1.501493
    (addr==142) ? 25193384 :   //   in=14.437500 val=1.501643
    (addr==143) ? 25195881 :   //   in=14.468750 val=1.501792
    (addr==144) ? 25198369 :   //   in=14.500000 val=1.501940
    (addr==145) ? 25200845 :   //   in=14.531250 val=1.502087
    (addr==146) ? 25203311 :   //   in=14.562500 val=1.502234
    (addr==147) ? 25205766 :   //   in=14.593750 val=1.502381
    (addr==148) ? 25208211 :   //   in=14.625000 val=1.502527
    (addr==149) ? 25210646 :   //   in=14.656250 val=1.502672
    (addr==150) ? 25213070 :   //   in=14.687500 val=1.502816
    (addr==151) ? 25215484 :   //   in=14.718750 val=1.502960
    (addr==152) ? 25217888 :   //   in=14.750000 val=1.503103
    (addr==153) ? 25220282 :   //   in=14.781250 val=1.503246
    (addr==154) ? 25222666 :   //   in=14.812500 val=1.503388
    (addr==155) ? 25225039 :   //   in=14.843750 val=1.503530
    (addr==156) ? 25227403 :   //   in=14.875000 val=1.503670
    (addr==157) ? 25229757 :   //   in=14.906250 val=1.503811
    (addr==158) ? 25232101 :   //   in=14.937500 val=1.503950
    (addr==159) ? 25234436 :   //   in=14.968750 val=1.504090
    (addr==160) ? 25236760 :   //   in=15.000000 val=1.504228
    (addr==161) ? 25239075 :   //   in=15.031250 val=1.504366
    (addr==162) ? 25241381 :   //   in=15.062500 val=1.504504
    (addr==163) ? 25243677 :   //   in=15.093750 val=1.504640
    (addr==164) ? 25245963 :   //   in=15.125000 val=1.504777
    (addr==165) ? 25248241 :   //   in=15.156250 val=1.504912
    (addr==166) ? 25250508 :   //   in=15.187500 val=1.505048
    (addr==167) ? 25252767 :   //   in=15.218750 val=1.505182
    (addr==168) ? 25255016 :   //   in=15.250000 val=1.505316
    (addr==169) ? 25257256 :   //   in=15.281250 val=1.505450
    (addr==170) ? 25259487 :   //   in=15.312500 val=1.505583
    (addr==171) ? 25261710 :   //   in=15.343750 val=1.505715
    (addr==172) ? 25263923 :   //   in=15.375000 val=1.505847
    (addr==173) ? 25266127 :   //   in=15.406250 val=1.505979
    (addr==174) ? 25268322 :   //   in=15.437500 val=1.506109
    (addr==175) ? 25270508 :   //   in=15.468750 val=1.506240
    (addr==176) ? 25272686 :   //   in=15.500000 val=1.506369
    (addr==177) ? 25274855 :   //   in=15.531250 val=1.506499
    (addr==178) ? 25277015 :   //   in=15.562500 val=1.506628
    (addr==179) ? 25279166 :   //   in=15.593750 val=1.506756
    (addr==180) ? 25281309 :   //   in=15.625000 val=1.506883
    (addr==181) ? 25283444 :   //   in=15.656250 val=1.507011
    (addr==182) ? 25285570 :   //   in=15.687500 val=1.507137
    (addr==183) ? 25287687 :   //   in=15.718750 val=1.507264
    (addr==184) ? 25289797 :   //   in=15.750000 val=1.507389
    (addr==185) ? 25291898 :   //   in=15.781250 val=1.507515
    (addr==186) ? 25293990 :   //   in=15.812500 val=1.507639
    (addr==187) ? 25296075 :   //   in=15.843750 val=1.507764
    (addr==188) ? 25298151 :   //   in=15.875000 val=1.507887
    (addr==189) ? 25300219 :   //   in=15.906250 val=1.508011
    (addr==190) ? 25302279 :   //   in=15.937500 val=1.508133
    (addr==191) ? 25304331 :   //   in=15.968750 val=1.508256
    (addr==192) ? 25306375 :   //   in=16.000000 val=1.508378
    (addr==193) ? 25308411 :   //   in=16.031250 val=1.508499
    (addr==194) ? 25310439 :   //   in=16.062500 val=1.508620
    (addr==195) ? 25312459 :   //   in=16.093750 val=1.508740
    (addr==196) ? 25314472 :   //   in=16.125000 val=1.508860
    (addr==197) ? 25316477 :   //   in=16.156250 val=1.508980
    (addr==198) ? 25318474 :   //   in=16.187500 val=1.509099
    (addr==199) ? 25320463 :   //   in=16.218750 val=1.509217
    (addr==200) ? 25322445 :   //   in=16.250000 val=1.509335
    (addr==201) ? 25324419 :   //   in=16.281250 val=1.509453
    (addr==202) ? 25326386 :   //   in=16.312500 val=1.509570
    (addr==203) ? 25328345 :   //   in=16.343750 val=1.509687
    (addr==204) ? 25330297 :   //   in=16.375000 val=1.509803
    (addr==205) ? 25332241 :   //   in=16.406250 val=1.509919
    (addr==206) ? 25334178 :   //   in=16.437500 val=1.510035
    (addr==207) ? 25336108 :   //   in=16.468750 val=1.510150
    (addr==208) ? 25338030 :   //   in=16.500000 val=1.510264
    (addr==209) ? 25339945 :   //   in=16.531250 val=1.510378
    (addr==210) ? 25341853 :   //   in=16.562500 val=1.510492
    (addr==211) ? 25343754 :   //   in=16.593750 val=1.510605
    (addr==212) ? 25345647 :   //   in=16.625000 val=1.510718
    (addr==213) ? 25347534 :   //   in=16.656250 val=1.510831
    (addr==214) ? 25349413 :   //   in=16.687500 val=1.510943
    (addr==215) ? 25351286 :   //   in=16.718750 val=1.511054
    (addr==216) ? 25353151 :   //   in=16.750000 val=1.511166
    (addr==217) ? 25355010 :   //   in=16.781250 val=1.511276
    (addr==218) ? 25356862 :   //   in=16.812500 val=1.511387
    (addr==219) ? 25358707 :   //   in=16.843750 val=1.511497
    (addr==220) ? 25360545 :   //   in=16.875000 val=1.511606
    (addr==221) ? 25362376 :   //   in=16.906250 val=1.511715
    (addr==222) ? 25364201 :   //   in=16.937500 val=1.511824
    (addr==223) ? 25366018 :   //   in=16.968750 val=1.511933
    (addr==224) ? 25367830 :   //   in=17.000000 val=1.512041
    (addr==225) ? 25369634 :   //   in=17.031250 val=1.512148
    (addr==226) ? 25371432 :   //   in=17.062500 val=1.512255
    (addr==227) ? 25373224 :   //   in=17.093750 val=1.512362
    (addr==228) ? 25375009 :   //   in=17.125000 val=1.512468
    (addr==229) ? 25376787 :   //   in=17.156250 val=1.512574
    (addr==230) ? 25378559 :   //   in=17.187500 val=1.512680
    (addr==231) ? 25380325 :   //   in=17.218750 val=1.512785
    (addr==232) ? 25382084 :   //   in=17.250000 val=1.512890
    (addr==233) ? 25383837 :   //   in=17.281250 val=1.512995
    (addr==234) ? 25385583 :   //   in=17.312500 val=1.513099
    (addr==235) ? 25387324 :   //   in=17.343750 val=1.513202
    (addr==236) ? 25389058 :   //   in=17.375000 val=1.513306
    (addr==237) ? 25390786 :   //   in=17.406250 val=1.513409
    (addr==238) ? 25392507 :   //   in=17.437500 val=1.513511
    (addr==239) ? 25394223 :   //   in=17.468750 val=1.513614
    (addr==240) ? 25395932 :   //   in=17.500000 val=1.513716
    (addr==241) ? 25397636 :   //   in=17.531250 val=1.513817
    (addr==242) ? 25399333 :   //   in=17.562500 val=1.513918
    (addr==243) ? 25401024 :   //   in=17.593750 val=1.514019
    (addr==244) ? 25402709 :   //   in=17.625000 val=1.514120
    (addr==245) ? 25404389 :   //   in=17.656250 val=1.514220
    (addr==246) ? 25406062 :   //   in=17.687500 val=1.514319
    (addr==247) ? 25407730 :   //   in=17.718750 val=1.514419
    (addr==248) ? 25409392 :   //   in=17.750000 val=1.514518
    (addr==249) ? 25411048 :   //   in=17.781250 val=1.514616
    (addr==250) ? 25412698 :   //   in=17.812500 val=1.514715
    (addr==251) ? 25414342 :   //   in=17.843750 val=1.514813
    (addr==252) ? 25415981 :   //   in=17.875000 val=1.514911
    (addr==253) ? 25417614 :   //   in=17.906250 val=1.515008
    (addr==254) ? 25419241 :   //   in=17.937500 val=1.515105
    (addr==255) ? 25420862 :   //   in=17.968750 val=1.515202
    (addr==256) ? 25422478 :   //   in=18.000000 val=1.515298
    (addr==257) ? 25424089 :   //   in=18.031250 val=1.515394
    (addr==258) ? 25425694 :   //   in=18.062500 val=1.515489
    (addr==259) ? 25427293 :   //   in=18.093750 val=1.515585
    (addr==260) ? 25428887 :   //   in=18.125000 val=1.515680
    (addr==261) ? 25430475 :   //   in=18.156250 val=1.515774
    (addr==262) ? 25432058 :   //   in=18.187500 val=1.515869
    (addr==263) ? 25433636 :   //   in=18.218750 val=1.515963
    (addr==264) ? 25435208 :   //   in=18.250000 val=1.516057
    (addr==265) ? 25436774 :   //   in=18.281250 val=1.516150
    (addr==266) ? 25438336 :   //   in=18.312500 val=1.516243
    (addr==267) ? 25439892 :   //   in=18.343750 val=1.516336
    (addr==268) ? 25441443 :   //   in=18.375000 val=1.516428
    (addr==269) ? 25442988 :   //   in=18.406250 val=1.516520
    (addr==270) ? 25444529 :   //   in=18.437500 val=1.516612
    (addr==271) ? 25446064 :   //   in=18.468750 val=1.516704
    (addr==272) ? 25447594 :   //   in=18.500000 val=1.516795
    (addr==273) ? 25449119 :   //   in=18.531250 val=1.516886
    (addr==274) ? 25450639 :   //   in=18.562500 val=1.516976
    (addr==275) ? 25452153 :   //   in=18.593750 val=1.517067
    (addr==276) ? 25453663 :   //   in=18.625000 val=1.517157
    (addr==277) ? 25455167 :   //   in=18.656250 val=1.517246
    (addr==278) ? 25456667 :   //   in=18.687500 val=1.517336
    (addr==279) ? 25458161 :   //   in=18.718750 val=1.517425
    (addr==280) ? 25459651 :   //   in=18.750000 val=1.517513
    (addr==281) ? 25461135 :   //   in=18.781250 val=1.517602
    (addr==282) ? 25462615 :   //   in=18.812500 val=1.517690
    (addr==283) ? 25464090 :   //   in=18.843750 val=1.517778
    (addr==284) ? 25465560 :   //   in=18.875000 val=1.517866
    (addr==285) ? 25467025 :   //   in=18.906250 val=1.517953
    (addr==286) ? 25468485 :   //   in=18.937500 val=1.518040
    (addr==287) ? 25469941 :   //   in=18.968750 val=1.518127
    (addr==288) ? 25471391 :   //   in=19.000000 val=1.518213
    (addr==289) ? 25472837 :   //   in=19.031250 val=1.518299
    (addr==290) ? 25474279 :   //   in=19.062500 val=1.518385
    (addr==291) ? 25475715 :   //   in=19.093750 val=1.518471
    (addr==292) ? 25477147 :   //   in=19.125000 val=1.518556
    (addr==293) ? 25478574 :   //   in=19.156250 val=1.518641
    (addr==294) ? 25479997 :   //   in=19.187500 val=1.518726
    (addr==295) ? 25481414 :   //   in=19.218750 val=1.518811
    (addr==296) ? 25482828 :   //   in=19.250000 val=1.518895
    (addr==297) ? 25484237 :   //   in=19.281250 val=1.518979
    (addr==298) ? 25485641 :   //   in=19.312500 val=1.519063
    (addr==299) ? 25487040 :   //   in=19.343750 val=1.519146
    (addr==300) ? 25488436 :   //   in=19.375000 val=1.519229
    (addr==301) ? 25489826 :   //   in=19.406250 val=1.519312
    (addr==302) ? 25491213 :   //   in=19.437500 val=1.519395
    (addr==303) ? 25492594 :   //   in=19.468750 val=1.519477
    (addr==304) ? 25493972 :   //   in=19.500000 val=1.519559
    (addr==305) ? 25495345 :   //   in=19.531250 val=1.519641
    (addr==306) ? 25496713 :   //   in=19.562500 val=1.519723
    (addr==307) ? 25498078 :   //   in=19.593750 val=1.519804
    (addr==308) ? 25499438 :   //   in=19.625000 val=1.519885
    (addr==309) ? 25500793 :   //   in=19.656250 val=1.519966
    (addr==310) ? 25502144 :   //   in=19.687500 val=1.520046
    (addr==311) ? 25503492 :   //   in=19.718750 val=1.520127
    (addr==312) ? 25504834 :   //   in=19.750000 val=1.520207
    (addr==313) ? 25506173 :   //   in=19.781250 val=1.520286
    (addr==314) ? 25507507 :   //   in=19.812500 val=1.520366
    (addr==315) ? 25508837 :   //   in=19.843750 val=1.520445
    (addr==316) ? 25510163 :   //   in=19.875000 val=1.520524
    (addr==317) ? 25511485 :   //   in=19.906250 val=1.520603
    (addr==318) ? 25512803 :   //   in=19.937500 val=1.520682
    (addr==319) ? 25514116 :   //   in=19.968750 val=1.520760
    (addr==320) ? 25515426 :   //   in=20.000000 val=1.520838
    (addr==321) ? 25516731 :   //   in=20.031250 val=1.520916
    (addr==322) ? 25518033 :   //   in=20.062500 val=1.520993
    (addr==323) ? 25519330 :   //   in=20.093750 val=1.521071
    (addr==324) ? 25520623 :   //   in=20.125000 val=1.521148
    (addr==325) ? 25521913 :   //   in=20.156250 val=1.521225
    (addr==326) ? 25523198 :   //   in=20.187500 val=1.521301
    (addr==327) ? 25524479 :   //   in=20.218750 val=1.521378
    (addr==328) ? 25525757 :   //   in=20.250000 val=1.521454
    (addr==329) ? 25527030 :   //   in=20.281250 val=1.521530
    (addr==330) ? 25528300 :   //   in=20.312500 val=1.521605
    (addr==331) ? 25529566 :   //   in=20.343750 val=1.521681
    (addr==332) ? 25530827 :   //   in=20.375000 val=1.521756
    (addr==333) ? 25532085 :   //   in=20.406250 val=1.521831
    (addr==334) ? 25533339 :   //   in=20.437500 val=1.521906
    (addr==335) ? 25534590 :   //   in=20.468750 val=1.521980
    (addr==336) ? 25535836 :   //   in=20.500000 val=1.522054
    (addr==337) ? 25537079 :   //   in=20.531250 val=1.522129
    (addr==338) ? 25538318 :   //   in=20.562500 val=1.522202
    (addr==339) ? 25539553 :   //   in=20.593750 val=1.522276
    (addr==340) ? 25540785 :   //   in=20.625000 val=1.522349
    (addr==341) ? 25542012 :   //   in=20.656250 val=1.522423
    (addr==342) ? 25543236 :   //   in=20.687500 val=1.522496
    (addr==343) ? 25544457 :   //   in=20.718750 val=1.522568
    (addr==344) ? 25545673 :   //   in=20.750000 val=1.522641
    (addr==345) ? 25546886 :   //   in=20.781250 val=1.522713
    (addr==346) ? 25548096 :   //   in=20.812500 val=1.522785
    (addr==347) ? 25549302 :   //   in=20.843750 val=1.522857
    (addr==348) ? 25550504 :   //   in=20.875000 val=1.522929
    (addr==349) ? 25551702 :   //   in=20.906250 val=1.523000
    (addr==350) ? 25552897 :   //   in=20.937500 val=1.523071
    (addr==351) ? 25554089 :   //   in=20.968750 val=1.523142
    (addr==352) ? 25555277 :   //   in=21.000000 val=1.523213
    (addr==353) ? 25556461 :   //   in=21.031250 val=1.523284
    (addr==354) ? 25557642 :   //   in=21.062500 val=1.523354
    (addr==355) ? 25558820 :   //   in=21.093750 val=1.523424
    (addr==356) ? 25559993 :   //   in=21.125000 val=1.523494
    (addr==357) ? 25561164 :   //   in=21.156250 val=1.523564
    (addr==358) ? 25562331 :   //   in=21.187500 val=1.523634
    (addr==359) ? 25563495 :   //   in=21.218750 val=1.523703
    (addr==360) ? 25564655 :   //   in=21.250000 val=1.523772
    (addr==361) ? 25565812 :   //   in=21.281250 val=1.523841
    (addr==362) ? 25566965 :   //   in=21.312500 val=1.523910
    (addr==363) ? 25568115 :   //   in=21.343750 val=1.523978
    (addr==364) ? 25569262 :   //   in=21.375000 val=1.524047
    (addr==365) ? 25570405 :   //   in=21.406250 val=1.524115
    (addr==366) ? 25571545 :   //   in=21.437500 val=1.524183
    (addr==367) ? 25572682 :   //   in=21.468750 val=1.524251
    (addr==368) ? 25573815 :   //   in=21.500000 val=1.524318
    (addr==369) ? 25574945 :   //   in=21.531250 val=1.524386
    (addr==370) ? 25576072 :   //   in=21.562500 val=1.524453
    (addr==371) ? 25577196 :   //   in=21.593750 val=1.524520
    (addr==372) ? 25578316 :   //   in=21.625000 val=1.524586
    (addr==373) ? 25579433 :   //   in=21.656250 val=1.524653
    (addr==374) ? 25580547 :   //   in=21.687500 val=1.524719
    (addr==375) ? 25581658 :   //   in=21.718750 val=1.524786
    (addr==376) ? 25582765 :   //   in=21.750000 val=1.524852
    (addr==377) ? 25583870 :   //   in=21.781250 val=1.524917
    (addr==378) ? 25584971 :   //   in=21.812500 val=1.524983
    (addr==379) ? 25586069 :   //   in=21.843750 val=1.525049
    (addr==380) ? 25587164 :   //   in=21.875000 val=1.525114
    (addr==381) ? 25588256 :   //   in=21.906250 val=1.525179
    (addr==382) ? 25589344 :   //   in=21.937500 val=1.525244
    (addr==383) ? 25590430 :   //   in=21.968750 val=1.525309
    (addr==384) ? 25591513 :   //   in=22.000000 val=1.525373
    (addr==385) ? 25592592 :   //   in=22.031250 val=1.525437
    (addr==386) ? 25593668 :   //   in=22.062500 val=1.525502
    (addr==387) ? 25594742 :   //   in=22.093750 val=1.525566
    (addr==388) ? 25595812 :   //   in=22.125000 val=1.525629
    (addr==389) ? 25596880 :   //   in=22.156250 val=1.525693
    (addr==390) ? 25597944 :   //   in=22.187500 val=1.525756
    (addr==391) ? 25599005 :   //   in=22.218750 val=1.525820
    (addr==392) ? 25600064 :   //   in=22.250000 val=1.525883
    (addr==393) ? 25601119 :   //   in=22.281250 val=1.525946
    (addr==394) ? 25602172 :   //   in=22.312500 val=1.526008
    (addr==395) ? 25603221 :   //   in=22.343750 val=1.526071
    (addr==396) ? 25604268 :   //   in=22.375000 val=1.526133
    (addr==397) ? 25605311 :   //   in=22.406250 val=1.526196
    (addr==398) ? 25606352 :   //   in=22.437500 val=1.526258
    (addr==399) ? 25607390 :   //   in=22.468750 val=1.526319
    (addr==400) ? 25608425 :   //   in=22.500000 val=1.526381
    (addr==401) ? 25609457 :   //   in=22.531250 val=1.526443
    (addr==402) ? 25610487 :   //   in=22.562500 val=1.526504
    (addr==403) ? 25611513 :   //   in=22.593750 val=1.526565
    (addr==404) ? 25612537 :   //   in=22.625000 val=1.526626
    (addr==405) ? 25613557 :   //   in=22.656250 val=1.526687
    (addr==406) ? 25614575 :   //   in=22.687500 val=1.526748
    (addr==407) ? 25615591 :   //   in=22.718750 val=1.526808
    (addr==408) ? 25616603 :   //   in=22.750000 val=1.526869
    (addr==409) ? 25617613 :   //   in=22.781250 val=1.526929
    (addr==410) ? 25618620 :   //   in=22.812500 val=1.526989
    (addr==411) ? 25619624 :   //   in=22.843750 val=1.527049
    (addr==412) ? 25620625 :   //   in=22.875000 val=1.527108
    (addr==413) ? 25621624 :   //   in=22.906250 val=1.527168
    (addr==414) ? 25622620 :   //   in=22.937500 val=1.527227
    (addr==415) ? 25623613 :   //   in=22.968750 val=1.527286
    (addr==416) ? 25624604 :   //   in=23.000000 val=1.527345
    (addr==417) ? 25625592 :   //   in=23.031250 val=1.527404
    (addr==418) ? 25626577 :   //   in=23.062500 val=1.527463
    (addr==419) ? 25627559 :   //   in=23.093750 val=1.527522
    (addr==420) ? 25628539 :   //   in=23.125000 val=1.527580
    (addr==421) ? 25629517 :   //   in=23.156250 val=1.527638
    (addr==422) ? 25630491 :   //   in=23.187500 val=1.527696
    (addr==423) ? 25631463 :   //   in=23.218750 val=1.527754
    (addr==424) ? 25632433 :   //   in=23.250000 val=1.527812
    (addr==425) ? 25633399 :   //   in=23.281250 val=1.527870
    (addr==426) ? 25634364 :   //   in=23.312500 val=1.527927
    (addr==427) ? 25635325 :   //   in=23.343750 val=1.527984
    (addr==428) ? 25636284 :   //   in=23.375000 val=1.528042
    (addr==429) ? 25637241 :   //   in=23.406250 val=1.528099
    (addr==430) ? 25638195 :   //   in=23.437500 val=1.528156
    (addr==431) ? 25639146 :   //   in=23.468750 val=1.528212
    (addr==432) ? 25640095 :   //   in=23.500000 val=1.528269
    (addr==433) ? 25641042 :   //   in=23.531250 val=1.528325
    (addr==434) ? 25641985 :   //   in=23.562500 val=1.528381
    (addr==435) ? 25642927 :   //   in=23.593750 val=1.528438
    (addr==436) ? 25643866 :   //   in=23.625000 val=1.528494
    (addr==437) ? 25644802 :   //   in=23.656250 val=1.528549
    (addr==438) ? 25645736 :   //   in=23.687500 val=1.528605
    (addr==439) ? 25646668 :   //   in=23.718750 val=1.528661
    (addr==440) ? 25647597 :   //   in=23.750000 val=1.528716
    (addr==441) ? 25648523 :   //   in=23.781250 val=1.528771
    (addr==442) ? 25649448 :   //   in=23.812500 val=1.528826
    (addr==443) ? 25650369 :   //   in=23.843750 val=1.528881
    (addr==444) ? 25651289 :   //   in=23.875000 val=1.528936
    (addr==445) ? 25652206 :   //   in=23.906250 val=1.528991
    (addr==446) ? 25653120 :   //   in=23.937500 val=1.529045
    (addr==447) ? 25654032 :   //   in=23.968750 val=1.529100
    (addr==448) ? 25654942 :   //   in=24.000000 val=1.529154
    (addr==449) ? 25655850 :   //   in=24.031250 val=1.529208
    (addr==450) ? 25656755 :   //   in=24.062500 val=1.529262
    (addr==451) ? 25657658 :   //   in=24.093750 val=1.529316
    (addr==452) ? 25658558 :   //   in=24.125000 val=1.529369
    (addr==453) ? 25659456 :   //   in=24.156250 val=1.529423
    (addr==454) ? 25660352 :   //   in=24.187500 val=1.529476
    (addr==455) ? 25661245 :   //   in=24.218750 val=1.529529
    (addr==456) ? 25662137 :   //   in=24.250000 val=1.529583
    (addr==457) ? 25663025 :   //   in=24.281250 val=1.529636
    (addr==458) ? 25663912 :   //   in=24.312500 val=1.529688
    (addr==459) ? 25664796 :   //   in=24.343750 val=1.529741
    (addr==460) ? 25665678 :   //   in=24.375000 val=1.529794
    (addr==461) ? 25666558 :   //   in=24.406250 val=1.529846
    (addr==462) ? 25667436 :   //   in=24.437500 val=1.529898
    (addr==463) ? 25668311 :   //   in=24.468750 val=1.529951
    (addr==464) ? 25669184 :   //   in=24.500000 val=1.530003
    (addr==465) ? 25670055 :   //   in=24.531250 val=1.530055
    (addr==466) ? 25670924 :   //   in=24.562500 val=1.530106
    (addr==467) ? 25671790 :   //   in=24.593750 val=1.530158
    (addr==468) ? 25672655 :   //   in=24.625000 val=1.530209
    (addr==469) ? 25673517 :   //   in=24.656250 val=1.530261
    (addr==470) ? 25674377 :   //   in=24.687500 val=1.530312
    (addr==471) ? 25675234 :   //   in=24.718750 val=1.530363
    (addr==472) ? 25676090 :   //   in=24.750000 val=1.530414
    (addr==473) ? 25676943 :   //   in=24.781250 val=1.530465
    (addr==474) ? 25677795 :   //   in=24.812500 val=1.530516
    (addr==475) ? 25678644 :   //   in=24.843750 val=1.530566
    (addr==476) ? 25679491 :   //   in=24.875000 val=1.530617
    (addr==477) ? 25680336 :   //   in=24.906250 val=1.530667
    (addr==478) ? 25681178 :   //   in=24.937500 val=1.530718
    (addr==479) ? 25682019 :   //   in=24.968750 val=1.530768
    (addr==480) ? 25682858 :   //   in=25.000000 val=1.530818
    (addr==481) ? 25683694 :   //   in=25.031250 val=1.530867
    (addr==482) ? 25684529 :   //   in=25.062500 val=1.530917
    (addr==483) ? 25685361 :   //   in=25.093750 val=1.530967
    (addr==484) ? 25686191 :   //   in=25.125000 val=1.531016
    (addr==485) ? 25687019 :   //   in=25.156250 val=1.531066
    (addr==486) ? 25687845 :   //   in=25.187500 val=1.531115
    (addr==487) ? 25688670 :   //   in=25.218750 val=1.531164
    (addr==488) ? 25689492 :   //   in=25.250000 val=1.531213
    (addr==489) ? 25690312 :   //   in=25.281250 val=1.531262
    (addr==490) ? 25691130 :   //   in=25.312500 val=1.531311
    (addr==491) ? 25691946 :   //   in=25.343750 val=1.531359
    (addr==492) ? 25692760 :   //   in=25.375000 val=1.531408
    (addr==493) ? 25693572 :   //   in=25.406250 val=1.531456
    (addr==494) ? 25694382 :   //   in=25.437500 val=1.531505
    (addr==495) ? 25695190 :   //   in=25.468750 val=1.531553
    (addr==496) ? 25695996 :   //   in=25.500000 val=1.531601
    (addr==497) ? 25696800 :   //   in=25.531250 val=1.531649
    (addr==498) ? 25697602 :   //   in=25.562500 val=1.531696
    (addr==499) ? 25698402 :   //   in=25.593750 val=1.531744
    (addr==500) ? 25699200 :   //   in=25.625000 val=1.531792
    (addr==501) ? 25699996 :   //   in=25.656250 val=1.531839
    (addr==502) ? 25700791 :   //   in=25.687500 val=1.531887
    (addr==503) ? 25701583 :   //   in=25.718750 val=1.531934
    (addr==504) ? 25702374 :   //   in=25.750000 val=1.531981
    (addr==505) ? 25703162 :   //   in=25.781250 val=1.532028
    (addr==506) ? 25703949 :   //   in=25.812500 val=1.532075
    (addr==507) ? 25704734 :   //   in=25.843750 val=1.532122
    (addr==508) ? 25705516 :   //   in=25.875000 val=1.532168
    (addr==509) ? 25706297 :   //   in=25.906250 val=1.532215
    (addr==510) ? 25707077 :   //   in=25.937500 val=1.532261
    (addr==511) ? 25707854 :   //   in=25.968750 val=1.532308
    (addr==512) ? 25708629 :   //   in=26.000000 val=1.532354
    (addr==513) ? 25709403 :   //   in=26.031250 val=1.532400
    (addr==514) ? 25710174 :   //   in=26.062500 val=1.532446
    (addr==515) ? 25710944 :   //   in=26.093750 val=1.532492
    (addr==516) ? 25711712 :   //   in=26.125000 val=1.532537
    (addr==517) ? 25712478 :   //   in=26.156250 val=1.532583
    (addr==518) ? 25713242 :   //   in=26.187500 val=1.532629
    (addr==519) ? 25714005 :   //   in=26.218750 val=1.532674
    (addr==520) ? 25714766 :   //   in=26.250000 val=1.532720
    (addr==521) ? 25715525 :   //   in=26.281250 val=1.532765
    (addr==522) ? 25716282 :   //   in=26.312500 val=1.532810
    (addr==523) ? 25717037 :   //   in=26.343750 val=1.532855
    (addr==524) ? 25717790 :   //   in=26.375000 val=1.532900
    (addr==525) ? 25718542 :   //   in=26.406250 val=1.532945
    (addr==526) ? 25719292 :   //   in=26.437500 val=1.532989
    (addr==527) ? 25720040 :   //   in=26.468750 val=1.533034
    (addr==528) ? 25720787 :   //   in=26.500000 val=1.533078
    (addr==529) ? 25721531 :   //   in=26.531250 val=1.533123
    (addr==530) ? 25722274 :   //   in=26.562500 val=1.533167
    (addr==531) ? 25723015 :   //   in=26.593750 val=1.533211
    (addr==532) ? 25723755 :   //   in=26.625000 val=1.533255
    (addr==533) ? 25724492 :   //   in=26.656250 val=1.533299
    (addr==534) ? 25725228 :   //   in=26.687500 val=1.533343
    (addr==535) ? 25725963 :   //   in=26.718750 val=1.533387
    (addr==536) ? 25726695 :   //   in=26.750000 val=1.533431
    (addr==537) ? 25727426 :   //   in=26.781250 val=1.533474
    (addr==538) ? 25728155 :   //   in=26.812500 val=1.533518
    (addr==539) ? 25728882 :   //   in=26.843750 val=1.533561
    (addr==540) ? 25729608 :   //   in=26.875000 val=1.533604
    (addr==541) ? 25730332 :   //   in=26.906250 val=1.533647
    (addr==542) ? 25731055 :   //   in=26.937500 val=1.533690
    (addr==543) ? 25731775 :   //   in=26.968750 val=1.533733
    (addr==544) ? 25732494 :   //   in=27.000000 val=1.533776
    (addr==545) ? 25733212 :   //   in=27.031250 val=1.533819
    (addr==546) ? 25733927 :   //   in=27.062500 val=1.533862
    (addr==547) ? 25734641 :   //   in=27.093750 val=1.533904
    (addr==548) ? 25735354 :   //   in=27.125000 val=1.533947
    (addr==549) ? 25736065 :   //   in=27.156250 val=1.533989
    (addr==550) ? 25736774 :   //   in=27.187500 val=1.534031
    (addr==551) ? 25737481 :   //   in=27.218750 val=1.534073
    (addr==552) ? 25738187 :   //   in=27.250000 val=1.534116
    (addr==553) ? 25738892 :   //   in=27.281250 val=1.534158
    (addr==554) ? 25739594 :   //   in=27.312500 val=1.534199
    (addr==555) ? 25740295 :   //   in=27.343750 val=1.534241
    (addr==556) ? 25740995 :   //   in=27.375000 val=1.534283
    (addr==557) ? 25741693 :   //   in=27.406250 val=1.534324
    (addr==558) ? 25742389 :   //   in=27.437500 val=1.534366
    (addr==559) ? 25743084 :   //   in=27.468750 val=1.534407
    (addr==560) ? 25743777 :   //   in=27.500000 val=1.534449
    (addr==561) ? 25744468 :   //   in=27.531250 val=1.534490
    (addr==562) ? 25745158 :   //   in=27.562500 val=1.534531
    (addr==563) ? 25745847 :   //   in=27.593750 val=1.534572
    (addr==564) ? 25746534 :   //   in=27.625000 val=1.534613
    (addr==565) ? 25747219 :   //   in=27.656250 val=1.534654
    (addr==566) ? 25747903 :   //   in=27.687500 val=1.534695
    (addr==567) ? 25748585 :   //   in=27.718750 val=1.534735
    (addr==568) ? 25749266 :   //   in=27.750000 val=1.534776
    (addr==569) ? 25749945 :   //   in=27.781250 val=1.534816
    (addr==570) ? 25750623 :   //   in=27.812500 val=1.534857
    (addr==571) ? 25751299 :   //   in=27.843750 val=1.534897
    (addr==572) ? 25751974 :   //   in=27.875000 val=1.534937
    (addr==573) ? 25752647 :   //   in=27.906250 val=1.534977
    (addr==574) ? 25753318 :   //   in=27.937500 val=1.535017
    (addr==575) ? 25753988 :   //   in=27.968750 val=1.535057
    (addr==576) ? 25754657 :   //   in=28.000000 val=1.535097
    (addr==577) ? 25755324 :   //   in=28.031250 val=1.535137
    (addr==578) ? 25755990 :   //   in=28.062500 val=1.535177
    (addr==579) ? 25756654 :   //   in=28.093750 val=1.535216
    (addr==580) ? 25757317 :   //   in=28.125000 val=1.535256
    (addr==581) ? 25757978 :   //   in=28.156250 val=1.535295
    (addr==582) ? 25758638 :   //   in=28.187500 val=1.535334
    (addr==583) ? 25759296 :   //   in=28.218750 val=1.535374
    (addr==584) ? 25759953 :   //   in=28.250000 val=1.535413
    (addr==585) ? 25760608 :   //   in=28.281250 val=1.535452
    (addr==586) ? 25761262 :   //   in=28.312500 val=1.535491
    (addr==587) ? 25761915 :   //   in=28.343750 val=1.535530
    (addr==588) ? 25762566 :   //   in=28.375000 val=1.535569
    (addr==589) ? 25763216 :   //   in=28.406250 val=1.535607
    (addr==590) ? 25763864 :   //   in=28.437500 val=1.535646
    (addr==591) ? 25764511 :   //   in=28.468750 val=1.535685
    (addr==592) ? 25765156 :   //   in=28.500000 val=1.535723
    (addr==593) ? 25765800 :   //   in=28.531250 val=1.535761
    (addr==594) ? 25766442 :   //   in=28.562500 val=1.535800
    (addr==595) ? 25767084 :   //   in=28.593750 val=1.535838
    (addr==596) ? 25767723 :   //   in=28.625000 val=1.535876
    (addr==597) ? 25768362 :   //   in=28.656250 val=1.535914
    (addr==598) ? 25768999 :   //   in=28.687500 val=1.535952
    (addr==599) ? 25769634 :   //   in=28.718750 val=1.535990
    (addr==600) ? 25770269 :   //   in=28.750000 val=1.536028
    (addr==601) ? 25770901 :   //   in=28.781250 val=1.536065
    (addr==602) ? 25771533 :   //   in=28.812500 val=1.536103
    (addr==603) ? 25772163 :   //   in=28.843750 val=1.536141
    (addr==604) ? 25772792 :   //   in=28.875000 val=1.536178
    (addr==605) ? 25773419 :   //   in=28.906250 val=1.536216
    (addr==606) ? 25774045 :   //   in=28.937500 val=1.536253
    (addr==607) ? 25774670 :   //   in=28.968750 val=1.536290
    (addr==608) ? 25775293 :   //   in=29.000000 val=1.536327
    (addr==609) ? 25775915 :   //   in=29.031250 val=1.536364
    (addr==610) ? 25776536 :   //   in=29.062500 val=1.536401
    (addr==611) ? 25777155 :   //   in=29.093750 val=1.536438
    (addr==612) ? 25777773 :   //   in=29.125000 val=1.536475
    (addr==613) ? 25778390 :   //   in=29.156250 val=1.536512
    (addr==614) ? 25779005 :   //   in=29.187500 val=1.536548
    (addr==615) ? 25779619 :   //   in=29.218750 val=1.536585
    (addr==616) ? 25780232 :   //   in=29.250000 val=1.536622
    (addr==617) ? 25780843 :   //   in=29.281250 val=1.536658
    (addr==618) ? 25781454 :   //   in=29.312500 val=1.536694
    (addr==619) ? 25782062 :   //   in=29.343750 val=1.536731
    (addr==620) ? 25782670 :   //   in=29.375000 val=1.536767
    (addr==621) ? 25783276 :   //   in=29.406250 val=1.536803
    (addr==622) ? 25783881 :   //   in=29.437500 val=1.536839
    (addr==623) ? 25784485 :   //   in=29.468750 val=1.536875
    (addr==624) ? 25785087 :   //   in=29.500000 val=1.536911
    (addr==625) ? 25785688 :   //   in=29.531250 val=1.536947
    (addr==626) ? 25786288 :   //   in=29.562500 val=1.536983
    (addr==627) ? 25786887 :   //   in=29.593750 val=1.537018
    (addr==628) ? 25787484 :   //   in=29.625000 val=1.537054
    (addr==629) ? 25788080 :   //   in=29.656250 val=1.537089
    (addr==630) ? 25788675 :   //   in=29.687500 val=1.537125
    (addr==631) ? 25789269 :   //   in=29.718750 val=1.537160
    (addr==632) ? 25789861 :   //   in=29.750000 val=1.537196
    (addr==633) ? 25790452 :   //   in=29.781250 val=1.537231
    (addr==634) ? 25791042 :   //   in=29.812500 val=1.537266
    (addr==635) ? 25791631 :   //   in=29.843750 val=1.537301
    (addr==636) ? 25792218 :   //   in=29.875000 val=1.537336
    (addr==637) ? 25792804 :   //   in=29.906250 val=1.537371
    (addr==638) ? 25793389 :   //   in=29.937500 val=1.537406
    (addr==639) ? 25793973 :   //   in=29.968750 val=1.537441
    (addr==640) ? 25794555 :   //   in=30.000000 val=1.537475
    (addr==641) ? 25795137 :   //   in=30.031250 val=1.537510
    (addr==642) ? 25795717 :   //   in=30.062500 val=1.537545
    (addr==643) ? 25796295 :   //   in=30.093750 val=1.537579
    (addr==644) ? 25796873 :   //   in=30.125000 val=1.537613
    (addr==645) ? 25797450 :   //   in=30.156250 val=1.537648
    (addr==646) ? 25798025 :   //   in=30.187500 val=1.537682
    (addr==647) ? 25798599 :   //   in=30.218750 val=1.537716
    (addr==648) ? 25799172 :   //   in=30.250000 val=1.537751
    (addr==649) ? 25799744 :   //   in=30.281250 val=1.537785
    (addr==650) ? 25800314 :   //   in=30.312500 val=1.537819
    (addr==651) ? 25800884 :   //   in=30.343750 val=1.537853
    (addr==652) ? 25801452 :   //   in=30.375000 val=1.537886
    (addr==653) ? 25802019 :   //   in=30.406250 val=1.537920
    (addr==654) ? 25802585 :   //   in=30.437500 val=1.537954
    (addr==655) ? 25803150 :   //   in=30.468750 val=1.537988
    (addr==656) ? 25803713 :   //   in=30.500000 val=1.538021
    (addr==657) ? 25804276 :   //   in=30.531250 val=1.538055
    (addr==658) ? 25804837 :   //   in=30.562500 val=1.538088
    (addr==659) ? 25805397 :   //   in=30.593750 val=1.538122
    (addr==660) ? 25805956 :   //   in=30.625000 val=1.538155
    (addr==661) ? 25806514 :   //   in=30.656250 val=1.538188
    (addr==662) ? 25807070 :   //   in=30.687500 val=1.538221
    (addr==663) ? 25807626 :   //   in=30.718750 val=1.538254
    (addr==664) ? 25808180 :   //   in=30.750000 val=1.538287
    (addr==665) ? 25808734 :   //   in=30.781250 val=1.538320
    (addr==666) ? 25809286 :   //   in=30.812500 val=1.538353
    (addr==667) ? 25809837 :   //   in=30.843750 val=1.538386
    (addr==668) ? 25810387 :   //   in=30.875000 val=1.538419
    (addr==669) ? 25810936 :   //   in=30.906250 val=1.538452
    (addr==670) ? 25811484 :   //   in=30.937500 val=1.538484
    (addr==671) ? 25812030 :   //   in=30.968750 val=1.538517
    (addr==672) ? 25812576 :   //   in=31.000000 val=1.538549
    (addr==673) ? 25813120 :   //   in=31.031250 val=1.538582
    (addr==674) ? 25813664 :   //   in=31.062500 val=1.538614
    (addr==675) ? 25814206 :   //   in=31.093750 val=1.538647
    (addr==676) ? 25814747 :   //   in=31.125000 val=1.538679
    (addr==677) ? 25815287 :   //   in=31.156250 val=1.538711
    (addr==678) ? 25815826 :   //   in=31.187500 val=1.538743
    (addr==679) ? 25816364 :   //   in=31.218750 val=1.538775
    (addr==680) ? 25816901 :   //   in=31.250000 val=1.538807
    (addr==681) ? 25817437 :   //   in=31.281250 val=1.538839
    (addr==682) ? 25817971 :   //   in=31.312500 val=1.538871
    (addr==683) ? 25818505 :   //   in=31.343750 val=1.538903
    (addr==684) ? 25819038 :   //   in=31.375000 val=1.538935
    (addr==685) ? 25819569 :   //   in=31.406250 val=1.538966
    (addr==686) ? 25820100 :   //   in=31.437500 val=1.538998
    (addr==687) ? 25820629 :   //   in=31.468750 val=1.539029
    (addr==688) ? 25821158 :   //   in=31.500000 val=1.539061
    (addr==689) ? 25821685 :   //   in=31.531250 val=1.539092
    (addr==690) ? 25822211 :   //   in=31.562500 val=1.539124
    (addr==691) ? 25822736 :   //   in=31.593750 val=1.539155
    (addr==692) ? 25823261 :   //   in=31.625000 val=1.539186
    (addr==693) ? 25823784 :   //   in=31.656250 val=1.539217
    (addr==694) ? 25824306 :   //   in=31.687500 val=1.539249
    (addr==695) ? 25824827 :   //   in=31.718750 val=1.539280
    (addr==696) ? 25825347 :   //   in=31.750000 val=1.539311
    (addr==697) ? 25825866 :   //   in=31.781250 val=1.539342
    (addr==698) ? 25826384 :   //   in=31.812500 val=1.539372
    (addr==699) ? 25826901 :   //   in=31.843750 val=1.539403
    (addr==700) ? 25827417 :   //   in=31.875000 val=1.539434
    (addr==701) ? 25827932 :   //   in=31.906250 val=1.539465
    (addr==702) ? 25828446 :   //   in=31.937500 val=1.539495
    (addr==703) ? 25828959 :   //   in=31.968750 val=1.539526
    (addr==704) ? 25829471 :   //   in=32.000000 val=1.539556
    (addr==705) ? 25829982 :   //   in=32.031250 val=1.539587
    (addr==706) ? 25830492 :   //   in=32.062500 val=1.539617
    (addr==707) ? 25831001 :   //   in=32.093750 val=1.539648
    (addr==708) ? 25831509 :   //   in=32.125000 val=1.539678
    (addr==709) ? 25832016 :   //   in=32.156250 val=1.539708
    (addr==710) ? 25832522 :   //   in=32.187500 val=1.539738
    (addr==711) ? 25833028 :   //   in=32.218750 val=1.539768
    (addr==712) ? 25833532 :   //   in=32.250000 val=1.539799
    (addr==713) ? 25834035 :   //   in=32.281250 val=1.539828
    (addr==714) ? 25834537 :   //   in=32.312500 val=1.539858
    (addr==715) ? 25835038 :   //   in=32.343750 val=1.539888
    (addr==716) ? 25835538 :   //   in=32.375000 val=1.539918
    (addr==717) ? 25836038 :   //   in=32.406250 val=1.539948
    (addr==718) ? 25836536 :   //   in=32.437500 val=1.539978
    (addr==719) ? 25837033 :   //   in=32.468750 val=1.540007
    (addr==720) ? 25837530 :   //   in=32.500000 val=1.540037
    (addr==721) ? 25838025 :   //   in=32.531250 val=1.540066
    (addr==722) ? 25838519 :   //   in=32.562500 val=1.540096
    (addr==723) ? 25839013 :   //   in=32.593750 val=1.540125
    (addr==724) ? 25839506 :   //   in=32.625000 val=1.540155
    (addr==725) ? 25839997 :   //   in=32.656250 val=1.540184
    (addr==726) ? 25840488 :   //   in=32.687500 val=1.540213
    (addr==727) ? 25840978 :   //   in=32.718750 val=1.540242
    (addr==728) ? 25841466 :   //   in=32.750000 val=1.540271
    (addr==729) ? 25841954 :   //   in=32.781250 val=1.540301
    (addr==730) ? 25842441 :   //   in=32.812500 val=1.540330
    (addr==731) ? 25842927 :   //   in=32.843750 val=1.540359
    (addr==732) ? 25843413 :   //   in=32.875000 val=1.540387
    (addr==733) ? 25843897 :   //   in=32.906250 val=1.540416
    (addr==734) ? 25844380 :   //   in=32.937500 val=1.540445
    (addr==735) ? 25844862 :   //   in=32.968750 val=1.540474
    (addr==736) ? 25845344 :   //   in=33.000000 val=1.540503
    (addr==737) ? 25845824 :   //   in=33.031250 val=1.540531
    (addr==738) ? 25846304 :   //   in=33.062500 val=1.540560
    (addr==739) ? 25846783 :   //   in=33.093750 val=1.540588
    (addr==740) ? 25847261 :   //   in=33.125000 val=1.540617
    (addr==741) ? 25847737 :   //   in=33.156250 val=1.540645
    (addr==742) ? 25848214 :   //   in=33.187500 val=1.540674
    (addr==743) ? 25848689 :   //   in=33.218750 val=1.540702
    (addr==744) ? 25849163 :   //   in=33.250000 val=1.540730
    (addr==745) ? 25849636 :   //   in=33.281250 val=1.540758
    (addr==746) ? 25850109 :   //   in=33.312500 val=1.540787
    (addr==747) ? 25850580 :   //   in=33.343750 val=1.540815
    (addr==748) ? 25851051 :   //   in=33.375000 val=1.540843
    (addr==749) ? 25851521 :   //   in=33.406250 val=1.540871
    (addr==750) ? 25851990 :   //   in=33.437500 val=1.540899
    (addr==751) ? 25852458 :   //   in=33.468750 val=1.540927
    (addr==752) ? 25852925 :   //   in=33.500000 val=1.540954
    (addr==753) ? 25853391 :   //   in=33.531250 val=1.540982
    (addr==754) ? 25853857 :   //   in=33.562500 val=1.541010
    (addr==755) ? 25854321 :   //   in=33.593750 val=1.541038
    (addr==756) ? 25854785 :   //   in=33.625000 val=1.541065
    (addr==757) ? 25855248 :   //   in=33.656250 val=1.541093
    (addr==758) ? 25855710 :   //   in=33.687500 val=1.541120
    (addr==759) ? 25856171 :   //   in=33.718750 val=1.541148
    (addr==760) ? 25856631 :   //   in=33.750000 val=1.541175
    (addr==761) ? 25857091 :   //   in=33.781250 val=1.541203
    (addr==762) ? 25857550 :   //   in=33.812500 val=1.541230
    (addr==763) ? 25858007 :   //   in=33.843750 val=1.541257
    (addr==764) ? 25858464 :   //   in=33.875000 val=1.541285
    (addr==765) ? 25858920 :   //   in=33.906250 val=1.541312
    (addr==766) ? 25859375 :   //   in=33.937500 val=1.541339
    (addr==767) ? 25859830 :   //   in=33.968750 val=1.541366
    (addr==768) ? 25860283 :   //   in=34.000000 val=1.541393
    (addr==769) ? 25860736 :   //   in=34.031250 val=1.541420
    (addr==770) ? 25861188 :   //   in=34.062500 val=1.541447
    (addr==771) ? 25861639 :   //   in=34.093750 val=1.541474
    (addr==772) ? 25862089 :   //   in=34.125000 val=1.541501
    (addr==773) ? 25862539 :   //   in=34.156250 val=1.541527
    (addr==774) ? 25862987 :   //   in=34.187500 val=1.541554
    (addr==775) ? 25863435 :   //   in=34.218750 val=1.541581
    (addr==776) ? 25863882 :   //   in=34.250000 val=1.541608
    (addr==777) ? 25864328 :   //   in=34.281250 val=1.541634
    (addr==778) ? 25864774 :   //   in=34.312500 val=1.541661
    (addr==779) ? 25865218 :   //   in=34.343750 val=1.541687
    (addr==780) ? 25865662 :   //   in=34.375000 val=1.541714
    (addr==781) ? 25866105 :   //   in=34.406250 val=1.541740
    (addr==782) ? 25866547 :   //   in=34.437500 val=1.541766
    (addr==783) ? 25866988 :   //   in=34.468750 val=1.541793
    (addr==784) ? 25867429 :   //   in=34.500000 val=1.541819
    (addr==785) ? 25867868 :   //   in=34.531250 val=1.541845
    (addr==786) ? 25868307 :   //   in=34.562500 val=1.541871
    (addr==787) ? 25868746 :   //   in=34.593750 val=1.541897
    (addr==788) ? 25869183 :   //   in=34.625000 val=1.541923
    (addr==789) ? 25869619 :   //   in=34.656250 val=1.541950
    (addr==790) ? 25870055 :   //   in=34.687500 val=1.541975
    (addr==791) ? 25870490 :   //   in=34.718750 val=1.542001
    (addr==792) ? 25870924 :   //   in=34.750000 val=1.542027
    (addr==793) ? 25871358 :   //   in=34.781250 val=1.542053
    (addr==794) ? 25871790 :   //   in=34.812500 val=1.542079
    (addr==795) ? 25872222 :   //   in=34.843750 val=1.542105
    (addr==796) ? 25872653 :   //   in=34.875000 val=1.542130
    (addr==797) ? 25873084 :   //   in=34.906250 val=1.542156
    (addr==798) ? 25873513 :   //   in=34.937500 val=1.542182
    (addr==799) ? 25873942 :   //   in=34.968750 val=1.542207
    (addr==800) ? 25874370 :   //   in=35.000000 val=1.542233
    (addr==801) ? 25874797 :   //   in=35.031250 val=1.542258
    (addr==802) ? 25875224 :   //   in=35.062500 val=1.542284
    (addr==803) ? 25875650 :   //   in=35.093750 val=1.542309
    (addr==804) ? 25876075 :   //   in=35.125000 val=1.542334
    (addr==805) ? 25876499 :   //   in=35.156250 val=1.542360
    (addr==806) ? 25876922 :   //   in=35.187500 val=1.542385
    (addr==807) ? 25877345 :   //   in=35.218750 val=1.542410
    (addr==808) ? 25877767 :   //   in=35.250000 val=1.542435
    (addr==809) ? 25878188 :   //   in=35.281250 val=1.542460
    (addr==810) ? 25878609 :   //   in=35.312500 val=1.542485
    (addr==811) ? 25879028 :   //   in=35.343750 val=1.542510
    (addr==812) ? 25879447 :   //   in=35.375000 val=1.542535
    (addr==813) ? 25879866 :   //   in=35.406250 val=1.542560
    (addr==814) ? 25880283 :   //   in=35.437500 val=1.542585
    (addr==815) ? 25880700 :   //   in=35.468750 val=1.542610
    (addr==816) ? 25881116 :   //   in=35.500000 val=1.542635
    (addr==817) ? 25881531 :   //   in=35.531250 val=1.542660
    (addr==818) ? 25881946 :   //   in=35.562500 val=1.542684
    (addr==819) ? 25882360 :   //   in=35.593750 val=1.542709
    (addr==820) ? 25882773 :   //   in=35.625000 val=1.542734
    (addr==821) ? 25883185 :   //   in=35.656250 val=1.542758
    (addr==822) ? 25883597 :   //   in=35.687500 val=1.542783
    (addr==823) ? 25884008 :   //   in=35.718750 val=1.542807
    (addr==824) ? 25884418 :   //   in=35.750000 val=1.542832
    (addr==825) ? 25884828 :   //   in=35.781250 val=1.542856
    (addr==826) ? 25885237 :   //   in=35.812500 val=1.542880
    (addr==827) ? 25885645 :   //   in=35.843750 val=1.542905
    (addr==828) ? 25886052 :   //   in=35.875000 val=1.542929
    (addr==829) ? 25886459 :   //   in=35.906250 val=1.542953
    (addr==830) ? 25886865 :   //   in=35.937500 val=1.542977
    (addr==831) ? 25887270 :   //   in=35.968750 val=1.543002
    (addr==832) ? 25887675 :   //   in=36.000000 val=1.543026
    (addr==833) ? 25888079 :   //   in=36.031250 val=1.543050
    (addr==834) ? 25888482 :   //   in=36.062500 val=1.543074
    (addr==835) ? 25888884 :   //   in=36.093750 val=1.543098
    (addr==836) ? 25889286 :   //   in=36.125000 val=1.543122
    (addr==837) ? 25889687 :   //   in=36.156250 val=1.543146
    (addr==838) ? 25890088 :   //   in=36.187500 val=1.543170
    (addr==839) ? 25890487 :   //   in=36.218750 val=1.543193
    (addr==840) ? 25890886 :   //   in=36.250000 val=1.543217
    (addr==841) ? 25891285 :   //   in=36.281250 val=1.543241
    (addr==842) ? 25891682 :   //   in=36.312500 val=1.543265
    (addr==843) ? 25892079 :   //   in=36.343750 val=1.543288
    (addr==844) ? 25892476 :   //   in=36.375000 val=1.543312
    (addr==845) ? 25892871 :   //   in=36.406250 val=1.543335
    (addr==846) ? 25893266 :   //   in=36.437500 val=1.543359
    (addr==847) ? 25893660 :   //   in=36.468750 val=1.543382
    (addr==848) ? 25894054 :   //   in=36.500000 val=1.543406
    (addr==849) ? 25894447 :   //   in=36.531250 val=1.543429
    (addr==850) ? 25894839 :   //   in=36.562500 val=1.543453
    (addr==851) ? 25895231 :   //   in=36.593750 val=1.543476
    (addr==852) ? 25895622 :   //   in=36.625000 val=1.543499
    (addr==853) ? 25896012 :   //   in=36.656250 val=1.543523
    (addr==854) ? 25896401 :   //   in=36.687500 val=1.543546
    (addr==855) ? 25896790 :   //   in=36.718750 val=1.543569
    (addr==856) ? 25897179 :   //   in=36.750000 val=1.543592
    (addr==857) ? 25897566 :   //   in=36.781250 val=1.543615
    (addr==858) ? 25897953 :   //   in=36.812500 val=1.543638
    (addr==859) ? 25898339 :   //   in=36.843750 val=1.543661
    (addr==860) ? 25898725 :   //   in=36.875000 val=1.543684
    (addr==861) ? 25899110 :   //   in=36.906250 val=1.543707
    (addr==862) ? 25899494 :   //   in=36.937500 val=1.543730
    (addr==863) ? 25899878 :   //   in=36.968750 val=1.543753
    (addr==864) ? 25900261 :   //   in=37.000000 val=1.543776
    (addr==865) ? 25900643 :   //   in=37.031250 val=1.543799
    (addr==866) ? 25901025 :   //   in=37.062500 val=1.543821
    (addr==867) ? 25901406 :   //   in=37.093750 val=1.543844
    (addr==868) ? 25901786 :   //   in=37.125000 val=1.543867
    (addr==869) ? 25902166 :   //   in=37.156250 val=1.543889
    (addr==870) ? 25902545 :   //   in=37.187500 val=1.543912
    (addr==871) ? 25902924 :   //   in=37.218750 val=1.543935
    (addr==872) ? 25903302 :   //   in=37.250000 val=1.543957
    (addr==873) ? 25903679 :   //   in=37.281250 val=1.543980
    (addr==874) ? 25904056 :   //   in=37.312500 val=1.544002
    (addr==875) ? 25904432 :   //   in=37.343750 val=1.544024
    (addr==876) ? 25904807 :   //   in=37.375000 val=1.544047
    (addr==877) ? 25905182 :   //   in=37.406250 val=1.544069
    (addr==878) ? 25905556 :   //   in=37.437500 val=1.544091
    (addr==879) ? 25905929 :   //   in=37.468750 val=1.544114
    (addr==880) ? 25906302 :   //   in=37.500000 val=1.544136
    (addr==881) ? 25906675 :   //   in=37.531250 val=1.544158
    (addr==882) ? 25907046 :   //   in=37.562500 val=1.544180
    (addr==883) ? 25907417 :   //   in=37.593750 val=1.544202
    (addr==884) ? 25907788 :   //   in=37.625000 val=1.544225
    (addr==885) ? 25908157 :   //   in=37.656250 val=1.544247
    (addr==886) ? 25908527 :   //   in=37.687500 val=1.544269
    (addr==887) ? 25908895 :   //   in=37.718750 val=1.544291
    (addr==888) ? 25909263 :   //   in=37.750000 val=1.544312
    (addr==889) ? 25909630 :   //   in=37.781250 val=1.544334
    (addr==890) ? 25909997 :   //   in=37.812500 val=1.544356
    (addr==891) ? 25910363 :   //   in=37.843750 val=1.544378
    (addr==892) ? 25910729 :   //   in=37.875000 val=1.544400
    (addr==893) ? 25911094 :   //   in=37.906250 val=1.544422
    (addr==894) ? 25911458 :   //   in=37.937500 val=1.544443
    (addr==895) ? 25911822 :   //   in=37.968750 val=1.544465
    (addr==896) ? 25912185 :   //   in=38.000000 val=1.544487
    (addr==897) ? 25912547 :   //   in=38.031250 val=1.544508
    (addr==898) ? 25912909 :   //   in=38.062500 val=1.544530
    (addr==899) ? 25913271 :   //   in=38.093750 val=1.544551
    (addr==900) ? 25913632 :   //   in=38.125000 val=1.544573
    (addr==901) ? 25913992 :   //   in=38.156250 val=1.544594
    (addr==902) ? 25914351 :   //   in=38.187500 val=1.544616
    (addr==903) ? 25914710 :   //   in=38.218750 val=1.544637
    (addr==904) ? 25915069 :   //   in=38.250000 val=1.544658
    (addr==905) ? 25915426 :   //   in=38.281250 val=1.544680
    (addr==906) ? 25915784 :   //   in=38.312500 val=1.544701
    (addr==907) ? 25916140 :   //   in=38.343750 val=1.544722
    (addr==908) ? 25916496 :   //   in=38.375000 val=1.544744
    (addr==909) ? 25916852 :   //   in=38.406250 val=1.544765
    (addr==910) ? 25917207 :   //   in=38.437500 val=1.544786
    (addr==911) ? 25917561 :   //   in=38.468750 val=1.544807
    (addr==912) ? 25917915 :   //   in=38.500000 val=1.544828
    (addr==913) ? 25918268 :   //   in=38.531250 val=1.544849
    (addr==914) ? 25918621 :   //   in=38.562500 val=1.544870
    (addr==915) ? 25918973 :   //   in=38.593750 val=1.544891
    (addr==916) ? 25919324 :   //   in=38.625000 val=1.544912
    (addr==917) ? 25919675 :   //   in=38.656250 val=1.544933
    (addr==918) ? 25920025 :   //   in=38.687500 val=1.544954
    (addr==919) ? 25920375 :   //   in=38.718750 val=1.544975
    (addr==920) ? 25920724 :   //   in=38.750000 val=1.544996
    (addr==921) ? 25921073 :   //   in=38.781250 val=1.545016
    (addr==922) ? 25921421 :   //   in=38.812500 val=1.545037
    (addr==923) ? 25921769 :   //   in=38.843750 val=1.545058
    (addr==924) ? 25922116 :   //   in=38.875000 val=1.545079
    (addr==925) ? 25922462 :   //   in=38.906250 val=1.545099
    (addr==926) ? 25922808 :   //   in=38.937500 val=1.545120
    (addr==927) ? 25923153 :   //   in=38.968750 val=1.545140
    (addr==928) ? 25923498 :   //   in=39.000000 val=1.545161
    (addr==929) ? 25923842 :   //   in=39.031250 val=1.545181
    (addr==930) ? 25924186 :   //   in=39.062500 val=1.545202
    (addr==931) ? 25924529 :   //   in=39.093750 val=1.545222
    (addr==932) ? 25924871 :   //   in=39.125000 val=1.545243
    (addr==933) ? 25925213 :   //   in=39.156250 val=1.545263
    (addr==934) ? 25925555 :   //   in=39.187500 val=1.545284
    (addr==935) ? 25925896 :   //   in=39.218750 val=1.545304
    (addr==936) ? 25926236 :   //   in=39.250000 val=1.545324
    (addr==937) ? 25926576 :   //   in=39.281250 val=1.545344
    (addr==938) ? 25926915 :   //   in=39.312500 val=1.545365
    (addr==939) ? 25927254 :   //   in=39.343750 val=1.545385
    (addr==940) ? 25927592 :   //   in=39.375000 val=1.545405
    (addr==941) ? 25927930 :   //   in=39.406250 val=1.545425
    (addr==942) ? 25928267 :   //   in=39.437500 val=1.545445
    (addr==943) ? 25928604 :   //   in=39.468750 val=1.545465
    (addr==944) ? 25928940 :   //   in=39.500000 val=1.545485
    (addr==945) ? 25929275 :   //   in=39.531250 val=1.545505
    (addr==946) ? 25929610 :   //   in=39.562500 val=1.545525
    (addr==947) ? 25929945 :   //   in=39.593750 val=1.545545
    (addr==948) ? 25930279 :   //   in=39.625000 val=1.545565
    (addr==949) ? 25930612 :   //   in=39.656250 val=1.545585
    (addr==950) ? 25930945 :   //   in=39.687500 val=1.545605
    (addr==951) ? 25931278 :   //   in=39.718750 val=1.545625
    (addr==952) ? 25931609 :   //   in=39.750000 val=1.545644
    (addr==953) ? 25931941 :   //   in=39.781250 val=1.545664
    (addr==954) ? 25932272 :   //   in=39.812500 val=1.545684
    (addr==955) ? 25932602 :   //   in=39.843750 val=1.545704
    (addr==956) ? 25932932 :   //   in=39.875000 val=1.545723
    (addr==957) ? 25933261 :   //   in=39.906250 val=1.545743
    (addr==958) ? 25933590 :   //   in=39.937500 val=1.545762
    (addr==959) ? 25933918 :   //   in=39.968750 val=1.545782
    (addr==960) ? 25934246 :   //   in=40.000000 val=1.545802
    (addr==961) ? 25934573 :   //   in=40.031250 val=1.545821
    (addr==962) ? 25934900 :   //   in=40.062500 val=1.545841
    (addr==963) ? 25935226 :   //   in=40.093750 val=1.545860
    (addr==964) ? 25935552 :   //   in=40.125000 val=1.545879
    (addr==965) ? 25935877 :   //   in=40.156250 val=1.545899
    (addr==966) ? 25936201 :   //   in=40.187500 val=1.545918
    (addr==967) ? 25936526 :   //   in=40.218750 val=1.545937
    (addr==968) ? 25936849 :   //   in=40.250000 val=1.545957
    (addr==969) ? 25937172 :   //   in=40.281250 val=1.545976
    (addr==970) ? 25937495 :   //   in=40.312500 val=1.545995
    (addr==971) ? 25937817 :   //   in=40.343750 val=1.546014
    (addr==972) ? 25938139 :   //   in=40.375000 val=1.546034
    (addr==973) ? 25938460 :   //   in=40.406250 val=1.546053
    (addr==974) ? 25938781 :   //   in=40.437500 val=1.546072
    (addr==975) ? 25939101 :   //   in=40.468750 val=1.546091
    (addr==976) ? 25939421 :   //   in=40.500000 val=1.546110
    (addr==977) ? 25939740 :   //   in=40.531250 val=1.546129
    (addr==978) ? 25940059 :   //   in=40.562500 val=1.546148
    (addr==979) ? 25940377 :   //   in=40.593750 val=1.546167
    (addr==980) ? 25940695 :   //   in=40.625000 val=1.546186
    (addr==981) ? 25941012 :   //   in=40.656250 val=1.546205
    (addr==982) ? 25941329 :   //   in=40.687500 val=1.546224
    (addr==983) ? 25941645 :   //   in=40.718750 val=1.546243
    (addr==984) ? 25941961 :   //   in=40.750000 val=1.546261
    (addr==985) ? 25942276 :   //   in=40.781250 val=1.546280
    (addr==986) ? 25942591 :   //   in=40.812500 val=1.546299
    (addr==987) ? 25942905 :   //   in=40.843750 val=1.546318
    (addr==988) ? 25943219 :   //   in=40.875000 val=1.546336
    (addr==989) ? 25943532 :   //   in=40.906250 val=1.546355
    (addr==990) ? 25943845 :   //   in=40.937500 val=1.546374
    (addr==991) ? 25944158 :   //   in=40.968750 val=1.546392
    (addr==992) ? 25944469 :   //   in=41.000000 val=1.546411
    (addr==993) ? 25944781 :   //   in=41.031250 val=1.546429
    (addr==994) ? 25945092 :   //   in=41.062500 val=1.546448
    (addr==995) ? 25945402 :   //   in=41.093750 val=1.546467
    (addr==996) ? 25945713 :   //   in=41.125000 val=1.546485
    (addr==997) ? 25946022 :   //   in=41.156250 val=1.546503
    (addr==998) ? 25946331 :   //   in=41.187500 val=1.546522
    (addr==999) ? 25946640 :   //   in=41.218750 val=1.546540
    (addr==1000) ? 25946948 :   //   in=41.250000 val=1.546559
    (addr==1001) ? 25947256 :   //   in=41.281250 val=1.546577
    (addr==1002) ? 25947563 :   //   in=41.312500 val=1.546595
    (addr==1003) ? 25947870 :   //   in=41.343750 val=1.546614
    (addr==1004) ? 25948176 :   //   in=41.375000 val=1.546632
    (addr==1005) ? 25948482 :   //   in=41.406250 val=1.546650
    (addr==1006) ? 25948787 :   //   in=41.437500 val=1.546668
    (addr==1007) ? 25949092 :   //   in=41.468750 val=1.546686
    (addr==1008) ? 25949397 :   //   in=41.500000 val=1.546705
    (addr==1009) ? 25949701 :   //   in=41.531250 val=1.546723
    (addr==1010) ? 25950004 :   //   in=41.562500 val=1.546741
    (addr==1011) ? 25950307 :   //   in=41.593750 val=1.546759
    (addr==1012) ? 25950610 :   //   in=41.625000 val=1.546777
    (addr==1013) ? 25950912 :   //   in=41.656250 val=1.546795
    (addr==1014) ? 25951214 :   //   in=41.687500 val=1.546813
    (addr==1015) ? 25951515 :   //   in=41.718750 val=1.546831
    (addr==1016) ? 25951816 :   //   in=41.750000 val=1.546849
    (addr==1017) ? 25952116 :   //   in=41.781250 val=1.546867
    (addr==1018) ? 25952416 :   //   in=41.812500 val=1.546885
    (addr==1019) ? 25952716 :   //   in=41.843750 val=1.546902
    (addr==1020) ? 25953015 :   //   in=41.875000 val=1.546920
    (addr==1021) ? 25953314 :   //   in=41.906250 val=1.546938
    (addr==1022) ? 25953612 :   //   in=41.937500 val=1.546956
    (addr==1023) ? 25953909 :   //   in=41.968750 val=1.546974
25'bx;
assign lastone = 25829471;
endmodule
