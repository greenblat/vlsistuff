`define NC100_RGF_BASEADDR    'h0
`define ADDR_REGA                                                'h0
`define ADDR_CONTROL0                                            'h4
`define ADDR_STATUSA                                             'h8
`define ADDR_REGB                                                'hc
`define ADDR_EXTERN                                              'h10
`define ADDR_ETH0TMP0                                            'h100
`define ADDR_ETH0TMP1                                            'h104
`define ADDR_ETH0TMP2                                            'h108
`define ADDR_ETH1TMP0                                            'h200
`define ADDR_ETH1TMP1                                            'h204
`define ADDR_ETH1TMP2                                            'h208
`define ADDR_ETH2TMP0                                            'h300
`define ADDR_ETH2TMP1                                            'h304
`define ADDR_ETH2TMP2                                            'h308
`define ADDR_ETH3TMP0                                            'h400
`define ADDR_ETH3TMP1                                            'h404
`define ADDR_ETH3TMP2                                            'h408
`define ADDR_WIDER                                               'h40c
`define ADDR_LONGER                                              'h41c
`define ADDR_RONLY                                               'h42c
`define ADDR_RONLY2                                              'h430
`define ADDR_LDST_RAM                                            'h800
