`celldefine
module INV (input A, output Y);
assign  Y = ! A;
endmodule
`endcelldefine
