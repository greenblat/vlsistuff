
    module x16 #(parameter IDWID=4, parameter DWID=64, parameter EXTRAS=8, parameter WSTRB=DWID/8) ( input clk, input rst_n

    ,output [IDWID-1:0] slv0_arid
    ,output [31:0] slv0_araddr
    ,output [7:0] slv0_arlen
    ,output [EXTRAS-1:0] slv0_arextras
    ,output [1:0] slv0_arburst
    ,output slv0_arvalid
    ,input slv0_arready
    ,input [IDWID-1:0] slv0_rid
    ,input [DWID-1:0] slv0_rdata
    ,input [1:0] slv0_rresp
    ,input slv0_rlast
    ,input slv0_rvalid
    ,output slv0_rready

    ,output [IDWID-1:0] slv0_awid
    ,output [31:0] slv0_awaddr
    ,output [7:0] slv0_awlen
    ,output [EXTRAS-1:0] slv0_awextras
    ,output [1:0] slv0_awburst
    ,output slv0_awvalid
    ,input slv0_awready
    ,output [DWID-1:0] slv0_wdata
    ,output [WSTRB-1:0] slv0_wstrb
    ,output slv0_wlast
    ,output slv0_wvalid
    ,input slv0_wready
    ,input [IDWID-1:0] slv0_bid
    ,input [1:0] slv0_bresp
    ,input slv0_bvalid
    ,output slv0_bready

    ,output [IDWID-1:0] slv1_arid
    ,output [31:0] slv1_araddr
    ,output [7:0] slv1_arlen
    ,output [EXTRAS-1:0] slv1_arextras
    ,output [1:0] slv1_arburst
    ,output slv1_arvalid
    ,input slv1_arready
    ,input [IDWID-1:0] slv1_rid
    ,input [DWID-1:0] slv1_rdata
    ,input [1:0] slv1_rresp
    ,input slv1_rlast
    ,input slv1_rvalid
    ,output slv1_rready

    ,output [IDWID-1:0] slv1_awid
    ,output [31:0] slv1_awaddr
    ,output [7:0] slv1_awlen
    ,output [EXTRAS-1:0] slv1_awextras
    ,output [1:0] slv1_awburst
    ,output slv1_awvalid
    ,input slv1_awready
    ,output [DWID-1:0] slv1_wdata
    ,output [WSTRB-1:0] slv1_wstrb
    ,output slv1_wlast
    ,output slv1_wvalid
    ,input slv1_wready
    ,input [IDWID-1:0] slv1_bid
    ,input [1:0] slv1_bresp
    ,input slv1_bvalid
    ,output slv1_bready

    ,output [IDWID-1:0] slv10_arid
    ,output [31:0] slv10_araddr
    ,output [7:0] slv10_arlen
    ,output [EXTRAS-1:0] slv10_arextras
    ,output [1:0] slv10_arburst
    ,output slv10_arvalid
    ,input slv10_arready
    ,input [IDWID-1:0] slv10_rid
    ,input [DWID-1:0] slv10_rdata
    ,input [1:0] slv10_rresp
    ,input slv10_rlast
    ,input slv10_rvalid
    ,output slv10_rready

    ,output [IDWID-1:0] slv10_awid
    ,output [31:0] slv10_awaddr
    ,output [7:0] slv10_awlen
    ,output [EXTRAS-1:0] slv10_awextras
    ,output [1:0] slv10_awburst
    ,output slv10_awvalid
    ,input slv10_awready
    ,output [DWID-1:0] slv10_wdata
    ,output [WSTRB-1:0] slv10_wstrb
    ,output slv10_wlast
    ,output slv10_wvalid
    ,input slv10_wready
    ,input [IDWID-1:0] slv10_bid
    ,input [1:0] slv10_bresp
    ,input slv10_bvalid
    ,output slv10_bready

    ,output [IDWID-1:0] slv11_arid
    ,output [31:0] slv11_araddr
    ,output [7:0] slv11_arlen
    ,output [EXTRAS-1:0] slv11_arextras
    ,output [1:0] slv11_arburst
    ,output slv11_arvalid
    ,input slv11_arready
    ,input [IDWID-1:0] slv11_rid
    ,input [DWID-1:0] slv11_rdata
    ,input [1:0] slv11_rresp
    ,input slv11_rlast
    ,input slv11_rvalid
    ,output slv11_rready

    ,output [IDWID-1:0] slv11_awid
    ,output [31:0] slv11_awaddr
    ,output [7:0] slv11_awlen
    ,output [EXTRAS-1:0] slv11_awextras
    ,output [1:0] slv11_awburst
    ,output slv11_awvalid
    ,input slv11_awready
    ,output [DWID-1:0] slv11_wdata
    ,output [WSTRB-1:0] slv11_wstrb
    ,output slv11_wlast
    ,output slv11_wvalid
    ,input slv11_wready
    ,input [IDWID-1:0] slv11_bid
    ,input [1:0] slv11_bresp
    ,input slv11_bvalid
    ,output slv11_bready

    ,output [IDWID-1:0] slv12_arid
    ,output [31:0] slv12_araddr
    ,output [7:0] slv12_arlen
    ,output [EXTRAS-1:0] slv12_arextras
    ,output [1:0] slv12_arburst
    ,output slv12_arvalid
    ,input slv12_arready
    ,input [IDWID-1:0] slv12_rid
    ,input [DWID-1:0] slv12_rdata
    ,input [1:0] slv12_rresp
    ,input slv12_rlast
    ,input slv12_rvalid
    ,output slv12_rready

    ,output [IDWID-1:0] slv12_awid
    ,output [31:0] slv12_awaddr
    ,output [7:0] slv12_awlen
    ,output [EXTRAS-1:0] slv12_awextras
    ,output [1:0] slv12_awburst
    ,output slv12_awvalid
    ,input slv12_awready
    ,output [DWID-1:0] slv12_wdata
    ,output [WSTRB-1:0] slv12_wstrb
    ,output slv12_wlast
    ,output slv12_wvalid
    ,input slv12_wready
    ,input [IDWID-1:0] slv12_bid
    ,input [1:0] slv12_bresp
    ,input slv12_bvalid
    ,output slv12_bready

    ,output [IDWID-1:0] slv13_arid
    ,output [31:0] slv13_araddr
    ,output [7:0] slv13_arlen
    ,output [EXTRAS-1:0] slv13_arextras
    ,output [1:0] slv13_arburst
    ,output slv13_arvalid
    ,input slv13_arready
    ,input [IDWID-1:0] slv13_rid
    ,input [DWID-1:0] slv13_rdata
    ,input [1:0] slv13_rresp
    ,input slv13_rlast
    ,input slv13_rvalid
    ,output slv13_rready

    ,output [IDWID-1:0] slv13_awid
    ,output [31:0] slv13_awaddr
    ,output [7:0] slv13_awlen
    ,output [EXTRAS-1:0] slv13_awextras
    ,output [1:0] slv13_awburst
    ,output slv13_awvalid
    ,input slv13_awready
    ,output [DWID-1:0] slv13_wdata
    ,output [WSTRB-1:0] slv13_wstrb
    ,output slv13_wlast
    ,output slv13_wvalid
    ,input slv13_wready
    ,input [IDWID-1:0] slv13_bid
    ,input [1:0] slv13_bresp
    ,input slv13_bvalid
    ,output slv13_bready

    ,output [IDWID-1:0] slv14_arid
    ,output [31:0] slv14_araddr
    ,output [7:0] slv14_arlen
    ,output [EXTRAS-1:0] slv14_arextras
    ,output [1:0] slv14_arburst
    ,output slv14_arvalid
    ,input slv14_arready
    ,input [IDWID-1:0] slv14_rid
    ,input [DWID-1:0] slv14_rdata
    ,input [1:0] slv14_rresp
    ,input slv14_rlast
    ,input slv14_rvalid
    ,output slv14_rready

    ,output [IDWID-1:0] slv14_awid
    ,output [31:0] slv14_awaddr
    ,output [7:0] slv14_awlen
    ,output [EXTRAS-1:0] slv14_awextras
    ,output [1:0] slv14_awburst
    ,output slv14_awvalid
    ,input slv14_awready
    ,output [DWID-1:0] slv14_wdata
    ,output [WSTRB-1:0] slv14_wstrb
    ,output slv14_wlast
    ,output slv14_wvalid
    ,input slv14_wready
    ,input [IDWID-1:0] slv14_bid
    ,input [1:0] slv14_bresp
    ,input slv14_bvalid
    ,output slv14_bready

    ,output [IDWID-1:0] slv15_arid
    ,output [31:0] slv15_araddr
    ,output [7:0] slv15_arlen
    ,output [EXTRAS-1:0] slv15_arextras
    ,output [1:0] slv15_arburst
    ,output slv15_arvalid
    ,input slv15_arready
    ,input [IDWID-1:0] slv15_rid
    ,input [DWID-1:0] slv15_rdata
    ,input [1:0] slv15_rresp
    ,input slv15_rlast
    ,input slv15_rvalid
    ,output slv15_rready

    ,output [IDWID-1:0] slv15_awid
    ,output [31:0] slv15_awaddr
    ,output [7:0] slv15_awlen
    ,output [EXTRAS-1:0] slv15_awextras
    ,output [1:0] slv15_awburst
    ,output slv15_awvalid
    ,input slv15_awready
    ,output [DWID-1:0] slv15_wdata
    ,output [WSTRB-1:0] slv15_wstrb
    ,output slv15_wlast
    ,output slv15_wvalid
    ,input slv15_wready
    ,input [IDWID-1:0] slv15_bid
    ,input [1:0] slv15_bresp
    ,input slv15_bvalid
    ,output slv15_bready

    ,output [IDWID-1:0] slv2_arid
    ,output [31:0] slv2_araddr
    ,output [7:0] slv2_arlen
    ,output [EXTRAS-1:0] slv2_arextras
    ,output [1:0] slv2_arburst
    ,output slv2_arvalid
    ,input slv2_arready
    ,input [IDWID-1:0] slv2_rid
    ,input [DWID-1:0] slv2_rdata
    ,input [1:0] slv2_rresp
    ,input slv2_rlast
    ,input slv2_rvalid
    ,output slv2_rready

    ,output [IDWID-1:0] slv2_awid
    ,output [31:0] slv2_awaddr
    ,output [7:0] slv2_awlen
    ,output [EXTRAS-1:0] slv2_awextras
    ,output [1:0] slv2_awburst
    ,output slv2_awvalid
    ,input slv2_awready
    ,output [DWID-1:0] slv2_wdata
    ,output [WSTRB-1:0] slv2_wstrb
    ,output slv2_wlast
    ,output slv2_wvalid
    ,input slv2_wready
    ,input [IDWID-1:0] slv2_bid
    ,input [1:0] slv2_bresp
    ,input slv2_bvalid
    ,output slv2_bready

    ,output [IDWID-1:0] slv3_arid
    ,output [31:0] slv3_araddr
    ,output [7:0] slv3_arlen
    ,output [EXTRAS-1:0] slv3_arextras
    ,output [1:0] slv3_arburst
    ,output slv3_arvalid
    ,input slv3_arready
    ,input [IDWID-1:0] slv3_rid
    ,input [DWID-1:0] slv3_rdata
    ,input [1:0] slv3_rresp
    ,input slv3_rlast
    ,input slv3_rvalid
    ,output slv3_rready

    ,output [IDWID-1:0] slv3_awid
    ,output [31:0] slv3_awaddr
    ,output [7:0] slv3_awlen
    ,output [EXTRAS-1:0] slv3_awextras
    ,output [1:0] slv3_awburst
    ,output slv3_awvalid
    ,input slv3_awready
    ,output [DWID-1:0] slv3_wdata
    ,output [WSTRB-1:0] slv3_wstrb
    ,output slv3_wlast
    ,output slv3_wvalid
    ,input slv3_wready
    ,input [IDWID-1:0] slv3_bid
    ,input [1:0] slv3_bresp
    ,input slv3_bvalid
    ,output slv3_bready

    ,output [IDWID-1:0] slv4_arid
    ,output [31:0] slv4_araddr
    ,output [7:0] slv4_arlen
    ,output [EXTRAS-1:0] slv4_arextras
    ,output [1:0] slv4_arburst
    ,output slv4_arvalid
    ,input slv4_arready
    ,input [IDWID-1:0] slv4_rid
    ,input [DWID-1:0] slv4_rdata
    ,input [1:0] slv4_rresp
    ,input slv4_rlast
    ,input slv4_rvalid
    ,output slv4_rready

    ,output [IDWID-1:0] slv4_awid
    ,output [31:0] slv4_awaddr
    ,output [7:0] slv4_awlen
    ,output [EXTRAS-1:0] slv4_awextras
    ,output [1:0] slv4_awburst
    ,output slv4_awvalid
    ,input slv4_awready
    ,output [DWID-1:0] slv4_wdata
    ,output [WSTRB-1:0] slv4_wstrb
    ,output slv4_wlast
    ,output slv4_wvalid
    ,input slv4_wready
    ,input [IDWID-1:0] slv4_bid
    ,input [1:0] slv4_bresp
    ,input slv4_bvalid
    ,output slv4_bready

    ,output [IDWID-1:0] slv5_arid
    ,output [31:0] slv5_araddr
    ,output [7:0] slv5_arlen
    ,output [EXTRAS-1:0] slv5_arextras
    ,output [1:0] slv5_arburst
    ,output slv5_arvalid
    ,input slv5_arready
    ,input [IDWID-1:0] slv5_rid
    ,input [DWID-1:0] slv5_rdata
    ,input [1:0] slv5_rresp
    ,input slv5_rlast
    ,input slv5_rvalid
    ,output slv5_rready

    ,output [IDWID-1:0] slv5_awid
    ,output [31:0] slv5_awaddr
    ,output [7:0] slv5_awlen
    ,output [EXTRAS-1:0] slv5_awextras
    ,output [1:0] slv5_awburst
    ,output slv5_awvalid
    ,input slv5_awready
    ,output [DWID-1:0] slv5_wdata
    ,output [WSTRB-1:0] slv5_wstrb
    ,output slv5_wlast
    ,output slv5_wvalid
    ,input slv5_wready
    ,input [IDWID-1:0] slv5_bid
    ,input [1:0] slv5_bresp
    ,input slv5_bvalid
    ,output slv5_bready

    ,output [IDWID-1:0] slv6_arid
    ,output [31:0] slv6_araddr
    ,output [7:0] slv6_arlen
    ,output [EXTRAS-1:0] slv6_arextras
    ,output [1:0] slv6_arburst
    ,output slv6_arvalid
    ,input slv6_arready
    ,input [IDWID-1:0] slv6_rid
    ,input [DWID-1:0] slv6_rdata
    ,input [1:0] slv6_rresp
    ,input slv6_rlast
    ,input slv6_rvalid
    ,output slv6_rready

    ,output [IDWID-1:0] slv6_awid
    ,output [31:0] slv6_awaddr
    ,output [7:0] slv6_awlen
    ,output [EXTRAS-1:0] slv6_awextras
    ,output [1:0] slv6_awburst
    ,output slv6_awvalid
    ,input slv6_awready
    ,output [DWID-1:0] slv6_wdata
    ,output [WSTRB-1:0] slv6_wstrb
    ,output slv6_wlast
    ,output slv6_wvalid
    ,input slv6_wready
    ,input [IDWID-1:0] slv6_bid
    ,input [1:0] slv6_bresp
    ,input slv6_bvalid
    ,output slv6_bready

    ,output [IDWID-1:0] slv7_arid
    ,output [31:0] slv7_araddr
    ,output [7:0] slv7_arlen
    ,output [EXTRAS-1:0] slv7_arextras
    ,output [1:0] slv7_arburst
    ,output slv7_arvalid
    ,input slv7_arready
    ,input [IDWID-1:0] slv7_rid
    ,input [DWID-1:0] slv7_rdata
    ,input [1:0] slv7_rresp
    ,input slv7_rlast
    ,input slv7_rvalid
    ,output slv7_rready

    ,output [IDWID-1:0] slv7_awid
    ,output [31:0] slv7_awaddr
    ,output [7:0] slv7_awlen
    ,output [EXTRAS-1:0] slv7_awextras
    ,output [1:0] slv7_awburst
    ,output slv7_awvalid
    ,input slv7_awready
    ,output [DWID-1:0] slv7_wdata
    ,output [WSTRB-1:0] slv7_wstrb
    ,output slv7_wlast
    ,output slv7_wvalid
    ,input slv7_wready
    ,input [IDWID-1:0] slv7_bid
    ,input [1:0] slv7_bresp
    ,input slv7_bvalid
    ,output slv7_bready

    ,output [IDWID-1:0] slv8_arid
    ,output [31:0] slv8_araddr
    ,output [7:0] slv8_arlen
    ,output [EXTRAS-1:0] slv8_arextras
    ,output [1:0] slv8_arburst
    ,output slv8_arvalid
    ,input slv8_arready
    ,input [IDWID-1:0] slv8_rid
    ,input [DWID-1:0] slv8_rdata
    ,input [1:0] slv8_rresp
    ,input slv8_rlast
    ,input slv8_rvalid
    ,output slv8_rready

    ,output [IDWID-1:0] slv8_awid
    ,output [31:0] slv8_awaddr
    ,output [7:0] slv8_awlen
    ,output [EXTRAS-1:0] slv8_awextras
    ,output [1:0] slv8_awburst
    ,output slv8_awvalid
    ,input slv8_awready
    ,output [DWID-1:0] slv8_wdata
    ,output [WSTRB-1:0] slv8_wstrb
    ,output slv8_wlast
    ,output slv8_wvalid
    ,input slv8_wready
    ,input [IDWID-1:0] slv8_bid
    ,input [1:0] slv8_bresp
    ,input slv8_bvalid
    ,output slv8_bready

    ,output [IDWID-1:0] slv9_arid
    ,output [31:0] slv9_araddr
    ,output [7:0] slv9_arlen
    ,output [EXTRAS-1:0] slv9_arextras
    ,output [1:0] slv9_arburst
    ,output slv9_arvalid
    ,input slv9_arready
    ,input [IDWID-1:0] slv9_rid
    ,input [DWID-1:0] slv9_rdata
    ,input [1:0] slv9_rresp
    ,input slv9_rlast
    ,input slv9_rvalid
    ,output slv9_rready

    ,output [IDWID-1:0] slv9_awid
    ,output [31:0] slv9_awaddr
    ,output [7:0] slv9_awlen
    ,output [EXTRAS-1:0] slv9_awextras
    ,output [1:0] slv9_awburst
    ,output slv9_awvalid
    ,input slv9_awready
    ,output [DWID-1:0] slv9_wdata
    ,output [WSTRB-1:0] slv9_wstrb
    ,output slv9_wlast
    ,output slv9_wvalid
    ,input slv9_wready
    ,input [IDWID-1:0] slv9_bid
    ,input [1:0] slv9_bresp
    ,input slv9_bvalid
    ,output slv9_bready

    ,input [IDWID-1:0] mst0_arid
    ,input [31:0] mst0_araddr
    ,input [7:0] mst0_arlen
    ,input [EXTRAS-1:0] mst0_arextras
    ,input [1:0] mst0_arburst
    ,input mst0_arvalid
    ,output mst0_arready
    ,output [IDWID-1:0] mst0_rid
    ,output [DWID-1:0] mst0_rdata
    ,output [1:0] mst0_rresp
    ,output mst0_rlast
    ,output mst0_rvalid
    ,input mst0_rready

    ,input [IDWID-1:0] mst0_awid
    ,input [31:0] mst0_awaddr
    ,input [7:0] mst0_awlen
    ,input [EXTRAS-1:0] mst0_awextras
    ,input [1:0] mst0_awburst
    ,input mst0_awvalid
    ,output mst0_awready
    ,input [DWID-1:0] mst0_wdata
    ,input [WSTRB-1:0] mst0_wstrb
    ,input mst0_wlast
    ,input mst0_wvalid
    ,output mst0_wready
    ,output [IDWID-1:0] mst0_bid
    ,output [1:0] mst0_bresp
    ,output mst0_bvalid
    ,input mst0_bready

    ,input [IDWID-1:0] mst1_arid
    ,input [31:0] mst1_araddr
    ,input [7:0] mst1_arlen
    ,input [EXTRAS-1:0] mst1_arextras
    ,input [1:0] mst1_arburst
    ,input mst1_arvalid
    ,output mst1_arready
    ,output [IDWID-1:0] mst1_rid
    ,output [DWID-1:0] mst1_rdata
    ,output [1:0] mst1_rresp
    ,output mst1_rlast
    ,output mst1_rvalid
    ,input mst1_rready

    ,input [IDWID-1:0] mst1_awid
    ,input [31:0] mst1_awaddr
    ,input [7:0] mst1_awlen
    ,input [EXTRAS-1:0] mst1_awextras
    ,input [1:0] mst1_awburst
    ,input mst1_awvalid
    ,output mst1_awready
    ,input [DWID-1:0] mst1_wdata
    ,input [WSTRB-1:0] mst1_wstrb
    ,input mst1_wlast
    ,input mst1_wvalid
    ,output mst1_wready
    ,output [IDWID-1:0] mst1_bid
    ,output [1:0] mst1_bresp
    ,output mst1_bvalid
    ,input mst1_bready

    ,input [IDWID-1:0] mst10_arid
    ,input [31:0] mst10_araddr
    ,input [7:0] mst10_arlen
    ,input [EXTRAS-1:0] mst10_arextras
    ,input [1:0] mst10_arburst
    ,input mst10_arvalid
    ,output mst10_arready
    ,output [IDWID-1:0] mst10_rid
    ,output [DWID-1:0] mst10_rdata
    ,output [1:0] mst10_rresp
    ,output mst10_rlast
    ,output mst10_rvalid
    ,input mst10_rready

    ,input [IDWID-1:0] mst10_awid
    ,input [31:0] mst10_awaddr
    ,input [7:0] mst10_awlen
    ,input [EXTRAS-1:0] mst10_awextras
    ,input [1:0] mst10_awburst
    ,input mst10_awvalid
    ,output mst10_awready
    ,input [DWID-1:0] mst10_wdata
    ,input [WSTRB-1:0] mst10_wstrb
    ,input mst10_wlast
    ,input mst10_wvalid
    ,output mst10_wready
    ,output [IDWID-1:0] mst10_bid
    ,output [1:0] mst10_bresp
    ,output mst10_bvalid
    ,input mst10_bready

    ,input [IDWID-1:0] mst11_arid
    ,input [31:0] mst11_araddr
    ,input [7:0] mst11_arlen
    ,input [EXTRAS-1:0] mst11_arextras
    ,input [1:0] mst11_arburst
    ,input mst11_arvalid
    ,output mst11_arready
    ,output [IDWID-1:0] mst11_rid
    ,output [DWID-1:0] mst11_rdata
    ,output [1:0] mst11_rresp
    ,output mst11_rlast
    ,output mst11_rvalid
    ,input mst11_rready

    ,input [IDWID-1:0] mst11_awid
    ,input [31:0] mst11_awaddr
    ,input [7:0] mst11_awlen
    ,input [EXTRAS-1:0] mst11_awextras
    ,input [1:0] mst11_awburst
    ,input mst11_awvalid
    ,output mst11_awready
    ,input [DWID-1:0] mst11_wdata
    ,input [WSTRB-1:0] mst11_wstrb
    ,input mst11_wlast
    ,input mst11_wvalid
    ,output mst11_wready
    ,output [IDWID-1:0] mst11_bid
    ,output [1:0] mst11_bresp
    ,output mst11_bvalid
    ,input mst11_bready

    ,input [IDWID-1:0] mst12_arid
    ,input [31:0] mst12_araddr
    ,input [7:0] mst12_arlen
    ,input [EXTRAS-1:0] mst12_arextras
    ,input [1:0] mst12_arburst
    ,input mst12_arvalid
    ,output mst12_arready
    ,output [IDWID-1:0] mst12_rid
    ,output [DWID-1:0] mst12_rdata
    ,output [1:0] mst12_rresp
    ,output mst12_rlast
    ,output mst12_rvalid
    ,input mst12_rready

    ,input [IDWID-1:0] mst12_awid
    ,input [31:0] mst12_awaddr
    ,input [7:0] mst12_awlen
    ,input [EXTRAS-1:0] mst12_awextras
    ,input [1:0] mst12_awburst
    ,input mst12_awvalid
    ,output mst12_awready
    ,input [DWID-1:0] mst12_wdata
    ,input [WSTRB-1:0] mst12_wstrb
    ,input mst12_wlast
    ,input mst12_wvalid
    ,output mst12_wready
    ,output [IDWID-1:0] mst12_bid
    ,output [1:0] mst12_bresp
    ,output mst12_bvalid
    ,input mst12_bready

    ,input [IDWID-1:0] mst13_arid
    ,input [31:0] mst13_araddr
    ,input [7:0] mst13_arlen
    ,input [EXTRAS-1:0] mst13_arextras
    ,input [1:0] mst13_arburst
    ,input mst13_arvalid
    ,output mst13_arready
    ,output [IDWID-1:0] mst13_rid
    ,output [DWID-1:0] mst13_rdata
    ,output [1:0] mst13_rresp
    ,output mst13_rlast
    ,output mst13_rvalid
    ,input mst13_rready

    ,input [IDWID-1:0] mst13_awid
    ,input [31:0] mst13_awaddr
    ,input [7:0] mst13_awlen
    ,input [EXTRAS-1:0] mst13_awextras
    ,input [1:0] mst13_awburst
    ,input mst13_awvalid
    ,output mst13_awready
    ,input [DWID-1:0] mst13_wdata
    ,input [WSTRB-1:0] mst13_wstrb
    ,input mst13_wlast
    ,input mst13_wvalid
    ,output mst13_wready
    ,output [IDWID-1:0] mst13_bid
    ,output [1:0] mst13_bresp
    ,output mst13_bvalid
    ,input mst13_bready

    ,input [IDWID-1:0] mst14_arid
    ,input [31:0] mst14_araddr
    ,input [7:0] mst14_arlen
    ,input [EXTRAS-1:0] mst14_arextras
    ,input [1:0] mst14_arburst
    ,input mst14_arvalid
    ,output mst14_arready
    ,output [IDWID-1:0] mst14_rid
    ,output [DWID-1:0] mst14_rdata
    ,output [1:0] mst14_rresp
    ,output mst14_rlast
    ,output mst14_rvalid
    ,input mst14_rready

    ,input [IDWID-1:0] mst14_awid
    ,input [31:0] mst14_awaddr
    ,input [7:0] mst14_awlen
    ,input [EXTRAS-1:0] mst14_awextras
    ,input [1:0] mst14_awburst
    ,input mst14_awvalid
    ,output mst14_awready
    ,input [DWID-1:0] mst14_wdata
    ,input [WSTRB-1:0] mst14_wstrb
    ,input mst14_wlast
    ,input mst14_wvalid
    ,output mst14_wready
    ,output [IDWID-1:0] mst14_bid
    ,output [1:0] mst14_bresp
    ,output mst14_bvalid
    ,input mst14_bready

    ,input [IDWID-1:0] mst15_arid
    ,input [31:0] mst15_araddr
    ,input [7:0] mst15_arlen
    ,input [EXTRAS-1:0] mst15_arextras
    ,input [1:0] mst15_arburst
    ,input mst15_arvalid
    ,output mst15_arready
    ,output [IDWID-1:0] mst15_rid
    ,output [DWID-1:0] mst15_rdata
    ,output [1:0] mst15_rresp
    ,output mst15_rlast
    ,output mst15_rvalid
    ,input mst15_rready

    ,input [IDWID-1:0] mst15_awid
    ,input [31:0] mst15_awaddr
    ,input [7:0] mst15_awlen
    ,input [EXTRAS-1:0] mst15_awextras
    ,input [1:0] mst15_awburst
    ,input mst15_awvalid
    ,output mst15_awready
    ,input [DWID-1:0] mst15_wdata
    ,input [WSTRB-1:0] mst15_wstrb
    ,input mst15_wlast
    ,input mst15_wvalid
    ,output mst15_wready
    ,output [IDWID-1:0] mst15_bid
    ,output [1:0] mst15_bresp
    ,output mst15_bvalid
    ,input mst15_bready

    ,input [IDWID-1:0] mst2_arid
    ,input [31:0] mst2_araddr
    ,input [7:0] mst2_arlen
    ,input [EXTRAS-1:0] mst2_arextras
    ,input [1:0] mst2_arburst
    ,input mst2_arvalid
    ,output mst2_arready
    ,output [IDWID-1:0] mst2_rid
    ,output [DWID-1:0] mst2_rdata
    ,output [1:0] mst2_rresp
    ,output mst2_rlast
    ,output mst2_rvalid
    ,input mst2_rready

    ,input [IDWID-1:0] mst2_awid
    ,input [31:0] mst2_awaddr
    ,input [7:0] mst2_awlen
    ,input [EXTRAS-1:0] mst2_awextras
    ,input [1:0] mst2_awburst
    ,input mst2_awvalid
    ,output mst2_awready
    ,input [DWID-1:0] mst2_wdata
    ,input [WSTRB-1:0] mst2_wstrb
    ,input mst2_wlast
    ,input mst2_wvalid
    ,output mst2_wready
    ,output [IDWID-1:0] mst2_bid
    ,output [1:0] mst2_bresp
    ,output mst2_bvalid
    ,input mst2_bready

    ,input [IDWID-1:0] mst3_arid
    ,input [31:0] mst3_araddr
    ,input [7:0] mst3_arlen
    ,input [EXTRAS-1:0] mst3_arextras
    ,input [1:0] mst3_arburst
    ,input mst3_arvalid
    ,output mst3_arready
    ,output [IDWID-1:0] mst3_rid
    ,output [DWID-1:0] mst3_rdata
    ,output [1:0] mst3_rresp
    ,output mst3_rlast
    ,output mst3_rvalid
    ,input mst3_rready

    ,input [IDWID-1:0] mst3_awid
    ,input [31:0] mst3_awaddr
    ,input [7:0] mst3_awlen
    ,input [EXTRAS-1:0] mst3_awextras
    ,input [1:0] mst3_awburst
    ,input mst3_awvalid
    ,output mst3_awready
    ,input [DWID-1:0] mst3_wdata
    ,input [WSTRB-1:0] mst3_wstrb
    ,input mst3_wlast
    ,input mst3_wvalid
    ,output mst3_wready
    ,output [IDWID-1:0] mst3_bid
    ,output [1:0] mst3_bresp
    ,output mst3_bvalid
    ,input mst3_bready

    ,input [IDWID-1:0] mst4_arid
    ,input [31:0] mst4_araddr
    ,input [7:0] mst4_arlen
    ,input [EXTRAS-1:0] mst4_arextras
    ,input [1:0] mst4_arburst
    ,input mst4_arvalid
    ,output mst4_arready
    ,output [IDWID-1:0] mst4_rid
    ,output [DWID-1:0] mst4_rdata
    ,output [1:0] mst4_rresp
    ,output mst4_rlast
    ,output mst4_rvalid
    ,input mst4_rready

    ,input [IDWID-1:0] mst4_awid
    ,input [31:0] mst4_awaddr
    ,input [7:0] mst4_awlen
    ,input [EXTRAS-1:0] mst4_awextras
    ,input [1:0] mst4_awburst
    ,input mst4_awvalid
    ,output mst4_awready
    ,input [DWID-1:0] mst4_wdata
    ,input [WSTRB-1:0] mst4_wstrb
    ,input mst4_wlast
    ,input mst4_wvalid
    ,output mst4_wready
    ,output [IDWID-1:0] mst4_bid
    ,output [1:0] mst4_bresp
    ,output mst4_bvalid
    ,input mst4_bready

    ,input [IDWID-1:0] mst5_arid
    ,input [31:0] mst5_araddr
    ,input [7:0] mst5_arlen
    ,input [EXTRAS-1:0] mst5_arextras
    ,input [1:0] mst5_arburst
    ,input mst5_arvalid
    ,output mst5_arready
    ,output [IDWID-1:0] mst5_rid
    ,output [DWID-1:0] mst5_rdata
    ,output [1:0] mst5_rresp
    ,output mst5_rlast
    ,output mst5_rvalid
    ,input mst5_rready

    ,input [IDWID-1:0] mst5_awid
    ,input [31:0] mst5_awaddr
    ,input [7:0] mst5_awlen
    ,input [EXTRAS-1:0] mst5_awextras
    ,input [1:0] mst5_awburst
    ,input mst5_awvalid
    ,output mst5_awready
    ,input [DWID-1:0] mst5_wdata
    ,input [WSTRB-1:0] mst5_wstrb
    ,input mst5_wlast
    ,input mst5_wvalid
    ,output mst5_wready
    ,output [IDWID-1:0] mst5_bid
    ,output [1:0] mst5_bresp
    ,output mst5_bvalid
    ,input mst5_bready

    ,input [IDWID-1:0] mst6_arid
    ,input [31:0] mst6_araddr
    ,input [7:0] mst6_arlen
    ,input [EXTRAS-1:0] mst6_arextras
    ,input [1:0] mst6_arburst
    ,input mst6_arvalid
    ,output mst6_arready
    ,output [IDWID-1:0] mst6_rid
    ,output [DWID-1:0] mst6_rdata
    ,output [1:0] mst6_rresp
    ,output mst6_rlast
    ,output mst6_rvalid
    ,input mst6_rready

    ,input [IDWID-1:0] mst6_awid
    ,input [31:0] mst6_awaddr
    ,input [7:0] mst6_awlen
    ,input [EXTRAS-1:0] mst6_awextras
    ,input [1:0] mst6_awburst
    ,input mst6_awvalid
    ,output mst6_awready
    ,input [DWID-1:0] mst6_wdata
    ,input [WSTRB-1:0] mst6_wstrb
    ,input mst6_wlast
    ,input mst6_wvalid
    ,output mst6_wready
    ,output [IDWID-1:0] mst6_bid
    ,output [1:0] mst6_bresp
    ,output mst6_bvalid
    ,input mst6_bready

    ,input [IDWID-1:0] mst7_arid
    ,input [31:0] mst7_araddr
    ,input [7:0] mst7_arlen
    ,input [EXTRAS-1:0] mst7_arextras
    ,input [1:0] mst7_arburst
    ,input mst7_arvalid
    ,output mst7_arready
    ,output [IDWID-1:0] mst7_rid
    ,output [DWID-1:0] mst7_rdata
    ,output [1:0] mst7_rresp
    ,output mst7_rlast
    ,output mst7_rvalid
    ,input mst7_rready

    ,input [IDWID-1:0] mst7_awid
    ,input [31:0] mst7_awaddr
    ,input [7:0] mst7_awlen
    ,input [EXTRAS-1:0] mst7_awextras
    ,input [1:0] mst7_awburst
    ,input mst7_awvalid
    ,output mst7_awready
    ,input [DWID-1:0] mst7_wdata
    ,input [WSTRB-1:0] mst7_wstrb
    ,input mst7_wlast
    ,input mst7_wvalid
    ,output mst7_wready
    ,output [IDWID-1:0] mst7_bid
    ,output [1:0] mst7_bresp
    ,output mst7_bvalid
    ,input mst7_bready

    ,input [IDWID-1:0] mst8_arid
    ,input [31:0] mst8_araddr
    ,input [7:0] mst8_arlen
    ,input [EXTRAS-1:0] mst8_arextras
    ,input [1:0] mst8_arburst
    ,input mst8_arvalid
    ,output mst8_arready
    ,output [IDWID-1:0] mst8_rid
    ,output [DWID-1:0] mst8_rdata
    ,output [1:0] mst8_rresp
    ,output mst8_rlast
    ,output mst8_rvalid
    ,input mst8_rready

    ,input [IDWID-1:0] mst8_awid
    ,input [31:0] mst8_awaddr
    ,input [7:0] mst8_awlen
    ,input [EXTRAS-1:0] mst8_awextras
    ,input [1:0] mst8_awburst
    ,input mst8_awvalid
    ,output mst8_awready
    ,input [DWID-1:0] mst8_wdata
    ,input [WSTRB-1:0] mst8_wstrb
    ,input mst8_wlast
    ,input mst8_wvalid
    ,output mst8_wready
    ,output [IDWID-1:0] mst8_bid
    ,output [1:0] mst8_bresp
    ,output mst8_bvalid
    ,input mst8_bready

    ,input [IDWID-1:0] mst9_arid
    ,input [31:0] mst9_araddr
    ,input [7:0] mst9_arlen
    ,input [EXTRAS-1:0] mst9_arextras
    ,input [1:0] mst9_arburst
    ,input mst9_arvalid
    ,output mst9_arready
    ,output [IDWID-1:0] mst9_rid
    ,output [DWID-1:0] mst9_rdata
    ,output [1:0] mst9_rresp
    ,output mst9_rlast
    ,output mst9_rvalid
    ,input mst9_rready

    ,input [IDWID-1:0] mst9_awid
    ,input [31:0] mst9_awaddr
    ,input [7:0] mst9_awlen
    ,input [EXTRAS-1:0] mst9_awextras
    ,input [1:0] mst9_awburst
    ,input mst9_awvalid
    ,output mst9_awready
    ,input [DWID-1:0] mst9_wdata
    ,input [WSTRB-1:0] mst9_wstrb
    ,input mst9_wlast
    ,input mst9_wvalid
    ,output mst9_wready
    ,output [IDWID-1:0] mst9_bid
    ,output [1:0] mst9_bresp
    ,output mst9_bvalid
    ,input mst9_bready
);

wire [IDWID-1:0] split0_merge0_arid ;
wire [31:0] split0_merge0_araddr ;
wire [7:0] split0_merge0_arlen ;
wire [EXTRAS-1:0] split0_merge0_arextras ;
wire [1:0] split0_merge0_arburst ;
wire split0_merge0_arvalid ;
wire split0_merge0_arready ;
wire [IDWID-1:0] split0_merge0_rid ;
wire [DWID-1:0] split0_merge0_rdata ;
wire [1:0] split0_merge0_rresp ;
wire split0_merge0_rlast ;
wire split0_merge0_rvalid ;
wire split0_merge0_rready ;

wire [IDWID-1:0] split0_merge0_awid ;
wire [31:0] split0_merge0_awaddr ;
wire [7:0] split0_merge0_awlen ;
wire [EXTRAS-1:0] split0_merge0_awextras ;
wire [1:0] split0_merge0_awburst ;
wire split0_merge0_awvalid ;
wire split0_merge0_awready ;
wire [DWID-1:0] split0_merge0_wdata ;
wire [WSTRB-1:0] split0_merge0_wstrb ;
wire split0_merge0_wlast ;
wire split0_merge0_wvalid ;
wire split0_merge0_wready ;
wire [IDWID-1:0] split0_merge0_bid ;
wire [1:0] split0_merge0_bresp ;
wire split0_merge0_bvalid ;
wire split0_merge0_bready ;


wire [IDWID-1:0] split0_merge1_arid ;
wire [31:0] split0_merge1_araddr ;
wire [7:0] split0_merge1_arlen ;
wire [EXTRAS-1:0] split0_merge1_arextras ;
wire [1:0] split0_merge1_arburst ;
wire split0_merge1_arvalid ;
wire split0_merge1_arready ;
wire [IDWID-1:0] split0_merge1_rid ;
wire [DWID-1:0] split0_merge1_rdata ;
wire [1:0] split0_merge1_rresp ;
wire split0_merge1_rlast ;
wire split0_merge1_rvalid ;
wire split0_merge1_rready ;

wire [IDWID-1:0] split0_merge1_awid ;
wire [31:0] split0_merge1_awaddr ;
wire [7:0] split0_merge1_awlen ;
wire [EXTRAS-1:0] split0_merge1_awextras ;
wire [1:0] split0_merge1_awburst ;
wire split0_merge1_awvalid ;
wire split0_merge1_awready ;
wire [DWID-1:0] split0_merge1_wdata ;
wire [WSTRB-1:0] split0_merge1_wstrb ;
wire split0_merge1_wlast ;
wire split0_merge1_wvalid ;
wire split0_merge1_wready ;
wire [IDWID-1:0] split0_merge1_bid ;
wire [1:0] split0_merge1_bresp ;
wire split0_merge1_bvalid ;
wire split0_merge1_bready ;


wire [IDWID-1:0] split0_merge2_arid ;
wire [31:0] split0_merge2_araddr ;
wire [7:0] split0_merge2_arlen ;
wire [EXTRAS-1:0] split0_merge2_arextras ;
wire [1:0] split0_merge2_arburst ;
wire split0_merge2_arvalid ;
wire split0_merge2_arready ;
wire [IDWID-1:0] split0_merge2_rid ;
wire [DWID-1:0] split0_merge2_rdata ;
wire [1:0] split0_merge2_rresp ;
wire split0_merge2_rlast ;
wire split0_merge2_rvalid ;
wire split0_merge2_rready ;

wire [IDWID-1:0] split0_merge2_awid ;
wire [31:0] split0_merge2_awaddr ;
wire [7:0] split0_merge2_awlen ;
wire [EXTRAS-1:0] split0_merge2_awextras ;
wire [1:0] split0_merge2_awburst ;
wire split0_merge2_awvalid ;
wire split0_merge2_awready ;
wire [DWID-1:0] split0_merge2_wdata ;
wire [WSTRB-1:0] split0_merge2_wstrb ;
wire split0_merge2_wlast ;
wire split0_merge2_wvalid ;
wire split0_merge2_wready ;
wire [IDWID-1:0] split0_merge2_bid ;
wire [1:0] split0_merge2_bresp ;
wire split0_merge2_bvalid ;
wire split0_merge2_bready ;


wire [IDWID-1:0] split0_merge3_arid ;
wire [31:0] split0_merge3_araddr ;
wire [7:0] split0_merge3_arlen ;
wire [EXTRAS-1:0] split0_merge3_arextras ;
wire [1:0] split0_merge3_arburst ;
wire split0_merge3_arvalid ;
wire split0_merge3_arready ;
wire [IDWID-1:0] split0_merge3_rid ;
wire [DWID-1:0] split0_merge3_rdata ;
wire [1:0] split0_merge3_rresp ;
wire split0_merge3_rlast ;
wire split0_merge3_rvalid ;
wire split0_merge3_rready ;

wire [IDWID-1:0] split0_merge3_awid ;
wire [31:0] split0_merge3_awaddr ;
wire [7:0] split0_merge3_awlen ;
wire [EXTRAS-1:0] split0_merge3_awextras ;
wire [1:0] split0_merge3_awburst ;
wire split0_merge3_awvalid ;
wire split0_merge3_awready ;
wire [DWID-1:0] split0_merge3_wdata ;
wire [WSTRB-1:0] split0_merge3_wstrb ;
wire split0_merge3_wlast ;
wire split0_merge3_wvalid ;
wire split0_merge3_wready ;
wire [IDWID-1:0] split0_merge3_bid ;
wire [1:0] split0_merge3_bresp ;
wire split0_merge3_bvalid ;
wire split0_merge3_bready ;


axi_4_splitter split0 (
     .clk(clk) ,.rst_n(rst_n)

    ,.araddr(mst0_araddr[31:0])
    ,.arburst(mst0_arburst[1:0])
    ,.arextras(mst0_arextras[(EXTRAS - 1):0])
    ,.arid(mst0_arid[(IDWID - 1):0])
    ,.arlen(mst0_arlen[7:0])
    ,.arready(mst0_arready)
    ,.arvalid(mst0_arvalid)
    ,.awaddr(mst0_awaddr[31:0])
    ,.awburst(mst0_awburst[1:0])
    ,.awextras(mst0_awextras[(EXTRAS - 1):0])
    ,.awid(mst0_awid[3:0])
    ,.awlen(mst0_awlen[7:0])
    ,.awready(mst0_awready)
    ,.awvalid(mst0_awvalid)
    ,.bid(mst0_bid[(IDWID - 1):0])
    ,.bready(mst0_bready)
    ,.bresp(mst0_bresp[1:0])
    ,.bvalid(mst0_bvalid)
    ,.rdata(mst0_rdata[(DWID - 1):0])
    ,.rid(mst0_rid[(IDWID - 1):0])
    ,.rlast(mst0_rlast)
    ,.rready(mst0_rready)
    ,.rresp(mst0_rresp[1:0])
    ,.rvalid(mst0_rvalid)
    ,.wdata(mst0_wdata[(DWID - 1):0])
    ,.wlast(mst0_wlast)
    ,.wready(mst0_wready)
    ,.wstrb(mst0_wstrb[(WSTRB - 1):0])
    ,.wvalid(mst0_wvalid)

    ,.a_araddr(split0_merge0_araddr[31:0])
    ,.a_arburst(split0_merge0_arburst[1:0])
    ,.a_arextras(split0_merge0_arextras[(EXTRAS - 1):0])
    ,.a_arid(split0_merge0_arid[(IDWID - 1):0])
    ,.a_arlen(split0_merge0_arlen[7:0])
    ,.a_arready(split0_merge0_arready)
    ,.a_arvalid(split0_merge0_arvalid)
    ,.a_awaddr(split0_merge0_awaddr[31:0])
    ,.a_awburst(split0_merge0_awburst[1:0])
    ,.a_awextras(split0_merge0_awextras[(EXTRAS - 1):0])
    ,.a_awid(split0_merge0_awid[(IDWID - 1):0])
    ,.a_awlen(split0_merge0_awlen[7:0])
    ,.a_awready(split0_merge0_awready)
    ,.a_awvalid(split0_merge0_awvalid)
    ,.a_bid(split0_merge0_bid[(IDWID - 1):0])
    ,.a_bready(split0_merge0_bready)
    ,.a_bresp(split0_merge0_bresp[1:0])
    ,.a_bvalid(split0_merge0_bvalid)
    ,.a_rdata(split0_merge0_rdata[(DWID - 1):0])
    ,.a_rid(split0_merge0_rid[(IDWID - 1):0])
    ,.a_rlast(split0_merge0_rlast)
    ,.a_rready(split0_merge0_rready)
    ,.a_rresp(split0_merge0_rresp[1:0])
    ,.a_rvalid(split0_merge0_rvalid)
    ,.a_wdata(split0_merge0_wdata[(DWID - 1):0])
    ,.a_wlast(split0_merge0_wlast)
    ,.a_wready(split0_merge0_wready)
    ,.a_wstrb(split0_merge0_wstrb[(WSTRB - 1):0])
    ,.a_wvalid(split0_merge0_wvalid)
    ,.b_araddr(split0_merge1_araddr[31:0])
    ,.b_arburst(split0_merge1_arburst[1:0])
    ,.b_arextras(split0_merge1_arextras[(EXTRAS - 1):0])
    ,.b_arid(split0_merge1_arid[(IDWID - 1):0])
    ,.b_arlen(split0_merge1_arlen[7:0])
    ,.b_arready(split0_merge1_arready)
    ,.b_arvalid(split0_merge1_arvalid)
    ,.b_awaddr(split0_merge1_awaddr[31:0])
    ,.b_awburst(split0_merge1_awburst[1:0])
    ,.b_awextras(split0_merge1_awextras[(EXTRAS - 1):0])
    ,.b_awid(split0_merge1_awid[(IDWID - 1):0])
    ,.b_awlen(split0_merge1_awlen[7:0])
    ,.b_awready(split0_merge1_awready)
    ,.b_awvalid(split0_merge1_awvalid)
    ,.b_bid(split0_merge1_bid[(IDWID - 1):0])
    ,.b_bready(split0_merge1_bready)
    ,.b_bresp(split0_merge1_bresp[1:0])
    ,.b_bvalid(split0_merge1_bvalid)
    ,.b_rdata(split0_merge1_rdata[(DWID - 1):0])
    ,.b_rid(split0_merge1_rid[(IDWID - 1):0])
    ,.b_rlast(split0_merge1_rlast)
    ,.b_rready(split0_merge1_rready)
    ,.b_rresp(split0_merge1_rresp[1:0])
    ,.b_rvalid(split0_merge1_rvalid)
    ,.b_wdata(split0_merge1_wdata[(DWID - 1):0])
    ,.b_wlast(split0_merge1_wlast)
    ,.b_wready(split0_merge1_wready)
    ,.b_wstrb(split0_merge1_wstrb[(WSTRB - 1):0])
    ,.b_wvalid(split0_merge1_wvalid)
    ,.c_araddr(split0_merge2_araddr[31:0])
    ,.c_arburst(split0_merge2_arburst[1:0])
    ,.c_arextras(split0_merge2_arextras[(EXTRAS - 1):0])
    ,.c_arid(split0_merge2_arid[(IDWID - 1):0])
    ,.c_arlen(split0_merge2_arlen[7:0])
    ,.c_arready(split0_merge2_arready)
    ,.c_arvalid(split0_merge2_arvalid)
    ,.c_awaddr(split0_merge2_awaddr[31:0])
    ,.c_awburst(split0_merge2_awburst[1:0])
    ,.c_awextras(split0_merge2_awextras[(EXTRAS - 1):0])
    ,.c_awid(split0_merge2_awid[(IDWID - 1):0])
    ,.c_awlen(split0_merge2_awlen[7:0])
    ,.c_awready(split0_merge2_awready)
    ,.c_awvalid(split0_merge2_awvalid)
    ,.c_bid(split0_merge2_bid[(IDWID - 1):0])
    ,.c_bready(split0_merge2_bready)
    ,.c_bresp(split0_merge2_bresp[1:0])
    ,.c_bvalid(split0_merge2_bvalid)
    ,.c_rdata(split0_merge2_rdata[(DWID - 1):0])
    ,.c_rid(split0_merge2_rid[(IDWID - 1):0])
    ,.c_rlast(split0_merge2_rlast)
    ,.c_rready(split0_merge2_rready)
    ,.c_rresp(split0_merge2_rresp[1:0])
    ,.c_rvalid(split0_merge2_rvalid)
    ,.c_wdata(split0_merge2_wdata[(DWID - 1):0])
    ,.c_wlast(split0_merge2_wlast)
    ,.c_wready(split0_merge2_wready)
    ,.c_wstrb(split0_merge2_wstrb[(WSTRB - 1):0])
    ,.c_wvalid(split0_merge2_wvalid)
    ,.d_araddr(split0_merge3_araddr[31:0])
    ,.d_arburst(split0_merge3_arburst[1:0])
    ,.d_arextras(split0_merge3_arextras[(EXTRAS - 1):0])
    ,.d_arid(split0_merge3_arid[(IDWID - 1):0])
    ,.d_arlen(split0_merge3_arlen[7:0])
    ,.d_arready(split0_merge3_arready)
    ,.d_arvalid(split0_merge3_arvalid)
    ,.d_awaddr(split0_merge3_awaddr[31:0])
    ,.d_awburst(split0_merge3_awburst[1:0])
    ,.d_awextras(split0_merge3_awextras[(EXTRAS - 1):0])
    ,.d_awid(split0_merge3_awid[(IDWID - 1):0])
    ,.d_awlen(split0_merge3_awlen[7:0])
    ,.d_awready(split0_merge3_awready)
    ,.d_awvalid(split0_merge3_awvalid)
    ,.d_bid(split0_merge3_bid[(IDWID - 1):0])
    ,.d_bready(split0_merge3_bready)
    ,.d_bresp(split0_merge3_bresp[1:0])
    ,.d_bvalid(split0_merge3_bvalid)
    ,.d_rdata(split0_merge3_rdata[(DWID - 1):0])
    ,.d_rid(split0_merge3_rid[(IDWID - 1):0])
    ,.d_rlast(split0_merge3_rlast)
    ,.d_rready(split0_merge3_rready)
    ,.d_rresp(split0_merge3_rresp[1:0])
    ,.d_rvalid(split0_merge3_rvalid)
    ,.d_wdata(split0_merge3_wdata[(DWID - 1):0])
    ,.d_wlast(split0_merge3_wlast)
    ,.d_wready(split0_merge3_wready)
    ,.d_wstrb(split0_merge3_wstrb[(WSTRB - 1):0])
    ,.d_wvalid(split0_merge3_wvalid)

);

wire [IDWID-1:0] merge0_split100_arid ;
wire [31:0] merge0_split100_araddr ;
wire [7:0] merge0_split100_arlen ;
wire [EXTRAS-1:0] merge0_split100_arextras ;
wire [1:0] merge0_split100_arburst ;
wire merge0_split100_arvalid ;
wire merge0_split100_arready ;
wire [IDWID-1:0] merge0_split100_rid ;
wire [DWID-1:0] merge0_split100_rdata ;
wire [1:0] merge0_split100_rresp ;
wire merge0_split100_rlast ;
wire merge0_split100_rvalid ;
wire merge0_split100_rready ;

wire [IDWID-1:0] merge0_split100_awid ;
wire [31:0] merge0_split100_awaddr ;
wire [7:0] merge0_split100_awlen ;
wire [EXTRAS-1:0] merge0_split100_awextras ;
wire [1:0] merge0_split100_awburst ;
wire merge0_split100_awvalid ;
wire merge0_split100_awready ;
wire [DWID-1:0] merge0_split100_wdata ;
wire [WSTRB-1:0] merge0_split100_wstrb ;
wire merge0_split100_wlast ;
wire merge0_split100_wvalid ;
wire merge0_split100_wready ;
wire [IDWID-1:0] merge0_split100_bid ;
wire [1:0] merge0_split100_bresp ;
wire merge0_split100_bvalid ;
wire merge0_split100_bready ;


wire [IDWID-1:0] split1_merge0_arid ;
wire [31:0] split1_merge0_araddr ;
wire [7:0] split1_merge0_arlen ;
wire [EXTRAS-1:0] split1_merge0_arextras ;
wire [1:0] split1_merge0_arburst ;
wire split1_merge0_arvalid ;
wire split1_merge0_arready ;
wire [IDWID-1:0] split1_merge0_rid ;
wire [DWID-1:0] split1_merge0_rdata ;
wire [1:0] split1_merge0_rresp ;
wire split1_merge0_rlast ;
wire split1_merge0_rvalid ;
wire split1_merge0_rready ;

wire [IDWID-1:0] split1_merge0_awid ;
wire [31:0] split1_merge0_awaddr ;
wire [7:0] split1_merge0_awlen ;
wire [EXTRAS-1:0] split1_merge0_awextras ;
wire [1:0] split1_merge0_awburst ;
wire split1_merge0_awvalid ;
wire split1_merge0_awready ;
wire [DWID-1:0] split1_merge0_wdata ;
wire [WSTRB-1:0] split1_merge0_wstrb ;
wire split1_merge0_wlast ;
wire split1_merge0_wvalid ;
wire split1_merge0_wready ;
wire [IDWID-1:0] split1_merge0_bid ;
wire [1:0] split1_merge0_bresp ;
wire split1_merge0_bvalid ;
wire split1_merge0_bready ;


wire [IDWID-1:0] split2_merge0_arid ;
wire [31:0] split2_merge0_araddr ;
wire [7:0] split2_merge0_arlen ;
wire [EXTRAS-1:0] split2_merge0_arextras ;
wire [1:0] split2_merge0_arburst ;
wire split2_merge0_arvalid ;
wire split2_merge0_arready ;
wire [IDWID-1:0] split2_merge0_rid ;
wire [DWID-1:0] split2_merge0_rdata ;
wire [1:0] split2_merge0_rresp ;
wire split2_merge0_rlast ;
wire split2_merge0_rvalid ;
wire split2_merge0_rready ;

wire [IDWID-1:0] split2_merge0_awid ;
wire [31:0] split2_merge0_awaddr ;
wire [7:0] split2_merge0_awlen ;
wire [EXTRAS-1:0] split2_merge0_awextras ;
wire [1:0] split2_merge0_awburst ;
wire split2_merge0_awvalid ;
wire split2_merge0_awready ;
wire [DWID-1:0] split2_merge0_wdata ;
wire [WSTRB-1:0] split2_merge0_wstrb ;
wire split2_merge0_wlast ;
wire split2_merge0_wvalid ;
wire split2_merge0_wready ;
wire [IDWID-1:0] split2_merge0_bid ;
wire [1:0] split2_merge0_bresp ;
wire split2_merge0_bvalid ;
wire split2_merge0_bready ;


wire [IDWID-1:0] split3_merge0_arid ;
wire [31:0] split3_merge0_araddr ;
wire [7:0] split3_merge0_arlen ;
wire [EXTRAS-1:0] split3_merge0_arextras ;
wire [1:0] split3_merge0_arburst ;
wire split3_merge0_arvalid ;
wire split3_merge0_arready ;
wire [IDWID-1:0] split3_merge0_rid ;
wire [DWID-1:0] split3_merge0_rdata ;
wire [1:0] split3_merge0_rresp ;
wire split3_merge0_rlast ;
wire split3_merge0_rvalid ;
wire split3_merge0_rready ;

wire [IDWID-1:0] split3_merge0_awid ;
wire [31:0] split3_merge0_awaddr ;
wire [7:0] split3_merge0_awlen ;
wire [EXTRAS-1:0] split3_merge0_awextras ;
wire [1:0] split3_merge0_awburst ;
wire split3_merge0_awvalid ;
wire split3_merge0_awready ;
wire [DWID-1:0] split3_merge0_wdata ;
wire [WSTRB-1:0] split3_merge0_wstrb ;
wire split3_merge0_wlast ;
wire split3_merge0_wvalid ;
wire split3_merge0_wready ;
wire [IDWID-1:0] split3_merge0_bid ;
wire [1:0] split3_merge0_bresp ;
wire split3_merge0_bvalid ;
wire split3_merge0_bready ;


axi_4_merger merge0 (
     .clk(clk),.rst_n(rst_n)
    ,.araddr(merge0_split100_araddr[31:0])
    ,.arburst(merge0_split100_arburst[1:0])
    ,.arextras(merge0_split100_arextras[(EXTRAS - 1):0])
    ,.arid(merge0_split100_arid[(IDWID - 1):0])
    ,.arlen(merge0_split100_arlen[7:0])
    ,.arready(merge0_split100_arready)
    ,.arvalid(merge0_split100_arvalid)
    ,.awaddr(merge0_split100_awaddr[31:0])
    ,.awburst(merge0_split100_awburst[1:0])
    ,.awextras(merge0_split100_awextras[(EXTRAS - 1):0])
    ,.awid(merge0_split100_awid[3:0])
    ,.awlen(merge0_split100_awlen[7:0])
    ,.awready(merge0_split100_awready)
    ,.awvalid(merge0_split100_awvalid)
    ,.bid(merge0_split100_bid[(IDWID - 1):0])
    ,.bready(merge0_split100_bready)
    ,.bresp(merge0_split100_bresp[1:0])
    ,.bvalid(merge0_split100_bvalid)
    ,.rid(merge0_split100_rid[(IDWID - 1):0])
    ,.rlast(merge0_split100_rlast)
    ,.rready(merge0_split100_rready)
    ,.rresp(merge0_split100_rresp[1:0])
    ,.rvalid(merge0_split100_rvalid)
    ,.rdata(merge0_split100_rdata[(DWID - 1):0])
    ,.wdata(merge0_split100_wdata[(DWID - 1):0])
    ,.wlast(merge0_split100_wlast)
    ,.wready(merge0_split100_wready)
    ,.wstrb(merge0_split100_wstrb[(WSTRB - 1):0])
    ,.wvalid(merge0_split100_wvalid)


    ,.a_araddr(split0_merge0_araddr[31:0])
    ,.a_arburst(split0_merge0_arburst[1:0])
    ,.a_arextras(split0_merge0_arextras[(EXTRAS - 1):0])
    ,.a_arid(split0_merge0_arid[(IDWID - 1):0])
    ,.a_arlen(split0_merge0_arlen[7:0])
    ,.a_arready(split0_merge0_arready)
    ,.a_arvalid(split0_merge0_arvalid)
    ,.a_awaddr(split0_merge0_awaddr[31:0])
    ,.a_awburst(split0_merge0_awburst[1:0])
    ,.a_awextras(split0_merge0_awextras[(EXTRAS - 1):0])
    ,.a_awid(split0_merge0_awid[(IDWID - 1):0])
    ,.a_awlen(split0_merge0_awlen[7:0])
    ,.a_awready(split0_merge0_awready)
    ,.a_awvalid(split0_merge0_awvalid)
    ,.a_bid(split0_merge0_bid[(IDWID - 1):0])
    ,.a_bready(split0_merge0_bready)
    ,.a_bresp(split0_merge0_bresp[1:0])
    ,.a_bvalid(split0_merge0_bvalid)
    ,.a_rdata(split0_merge0_rdata[(DWID - 1):0])
    ,.a_rid(split0_merge0_rid[(IDWID - 1):0])
    ,.a_rlast(split0_merge0_rlast)
    ,.a_rready(split0_merge0_rready)
    ,.a_rresp(split0_merge0_rresp[1:0])
    ,.a_rvalid(split0_merge0_rvalid)
    ,.a_wdata(split0_merge0_wdata[(DWID - 1):0])
    ,.a_wlast(split0_merge0_wlast)
    ,.a_wready(split0_merge0_wready)
    ,.a_wstrb(split0_merge0_wstrb[(WSTRB - 1):0])
    ,.a_wvalid(split0_merge0_wvalid)

    ,.b_araddr(split1_merge0_araddr[31:0])
    ,.b_arburst(split1_merge0_arburst[1:0])
    ,.b_arextras(split1_merge0_arextras[(EXTRAS - 1):0])
    ,.b_arid(split1_merge0_arid[(IDWID - 1):0])
    ,.b_arlen(split1_merge0_arlen[7:0])
    ,.b_arready(split1_merge0_arready)
    ,.b_arvalid(split1_merge0_arvalid)
    ,.b_awaddr(split1_merge0_awaddr[31:0])
    ,.b_awburst(split1_merge0_awburst[1:0])
    ,.b_awextras(split1_merge0_awextras[(EXTRAS - 1):0])
    ,.b_awid(split1_merge0_awid[(IDWID - 1):0])
    ,.b_awlen(split1_merge0_awlen[7:0])
    ,.b_awready(split1_merge0_awready)
    ,.b_awvalid(split1_merge0_awvalid)
    ,.b_bid(split1_merge0_bid[(IDWID - 1):0])
    ,.b_bready(split1_merge0_bready)
    ,.b_bresp(split1_merge0_bresp[1:0])
    ,.b_bvalid(split1_merge0_bvalid)
    ,.b_rdata(split1_merge0_rdata[(DWID - 1):0])
    ,.b_rid(split1_merge0_rid[(IDWID - 1):0])
    ,.b_rlast(split1_merge0_rlast)
    ,.b_rready(split1_merge0_rready)
    ,.b_rresp(split1_merge0_rresp[1:0])
    ,.b_rvalid(split1_merge0_rvalid)
    ,.b_wdata(split1_merge0_wdata[(DWID - 1):0])
    ,.b_wlast(split1_merge0_wlast)
    ,.b_wready(split1_merge0_wready)
    ,.b_wstrb(split1_merge0_wstrb[(WSTRB - 1):0])
    ,.b_wvalid(split1_merge0_wvalid)

    ,.c_araddr(split2_merge0_araddr[31:0])
    ,.c_arburst(split2_merge0_arburst[1:0])
    ,.c_arextras(split2_merge0_arextras[(EXTRAS - 1):0])
    ,.c_arid(split2_merge0_arid[(IDWID - 1):0])
    ,.c_arlen(split2_merge0_arlen[7:0])
    ,.c_arready(split2_merge0_arready)
    ,.c_arvalid(split2_merge0_arvalid)
    ,.c_awaddr(split2_merge0_awaddr[31:0])
    ,.c_awburst(split2_merge0_awburst[1:0])
    ,.c_awextras(split2_merge0_awextras[(EXTRAS - 1):0])
    ,.c_awid(split2_merge0_awid[(IDWID - 1):0])
    ,.c_awlen(split2_merge0_awlen[7:0])
    ,.c_awready(split2_merge0_awready)
    ,.c_awvalid(split2_merge0_awvalid)
    ,.c_bid(split2_merge0_bid[(IDWID - 1):0])
    ,.c_bready(split2_merge0_bready)
    ,.c_bresp(split2_merge0_bresp[1:0])
    ,.c_bvalid(split2_merge0_bvalid)
    ,.c_rdata(split2_merge0_rdata[(DWID - 1):0])
    ,.c_rid(split2_merge0_rid[(IDWID - 1):0])
    ,.c_rlast(split2_merge0_rlast)
    ,.c_rready(split2_merge0_rready)
    ,.c_rresp(split2_merge0_rresp[1:0])
    ,.c_rvalid(split2_merge0_rvalid)
    ,.c_wdata(split2_merge0_wdata[(DWID - 1):0])
    ,.c_wlast(split2_merge0_wlast)
    ,.c_wready(split2_merge0_wready)
    ,.c_wstrb(split2_merge0_wstrb[(WSTRB - 1):0])
    ,.c_wvalid(split2_merge0_wvalid)

    ,.d_araddr(split3_merge0_araddr[31:0])
    ,.d_arburst(split3_merge0_arburst[1:0])
    ,.d_arextras(split3_merge0_arextras[(EXTRAS - 1):0])
    ,.d_arid(split3_merge0_arid[(IDWID - 1):0])
    ,.d_arlen(split3_merge0_arlen[7:0])
    ,.d_arready(split3_merge0_arready)
    ,.d_arvalid(split3_merge0_arvalid)
    ,.d_awaddr(split3_merge0_awaddr[31:0])
    ,.d_awburst(split3_merge0_awburst[1:0])
    ,.d_awextras(split3_merge0_awextras[(EXTRAS - 1):0])
    ,.d_awid(split3_merge0_awid[(IDWID - 1):0])
    ,.d_awlen(split3_merge0_awlen[7:0])
    ,.d_awready(split3_merge0_awready)
    ,.d_awvalid(split3_merge0_awvalid)
    ,.d_bid(split3_merge0_bid[(IDWID - 1):0])
    ,.d_bready(split3_merge0_bready)
    ,.d_bresp(split3_merge0_bresp[1:0])
    ,.d_bvalid(split3_merge0_bvalid)
    ,.d_rdata(split3_merge0_rdata[(DWID - 1):0])
    ,.d_rid(split3_merge0_rid[(IDWID - 1):0])
    ,.d_rlast(split3_merge0_rlast)
    ,.d_rready(split3_merge0_rready)
    ,.d_rresp(split3_merge0_rresp[1:0])
    ,.d_rvalid(split3_merge0_rvalid)
    ,.d_wdata(split3_merge0_wdata[(DWID - 1):0])
    ,.d_wlast(split3_merge0_wlast)
    ,.d_wready(split3_merge0_wready)
    ,.d_wstrb(split3_merge0_wstrb[(WSTRB - 1):0])
    ,.d_wvalid(split3_merge0_wvalid)
);


wire [IDWID-1:0] merge1_split101_arid ;
wire [31:0] merge1_split101_araddr ;
wire [7:0] merge1_split101_arlen ;
wire [EXTRAS-1:0] merge1_split101_arextras ;
wire [1:0] merge1_split101_arburst ;
wire merge1_split101_arvalid ;
wire merge1_split101_arready ;
wire [IDWID-1:0] merge1_split101_rid ;
wire [DWID-1:0] merge1_split101_rdata ;
wire [1:0] merge1_split101_rresp ;
wire merge1_split101_rlast ;
wire merge1_split101_rvalid ;
wire merge1_split101_rready ;

wire [IDWID-1:0] merge1_split101_awid ;
wire [31:0] merge1_split101_awaddr ;
wire [7:0] merge1_split101_awlen ;
wire [EXTRAS-1:0] merge1_split101_awextras ;
wire [1:0] merge1_split101_awburst ;
wire merge1_split101_awvalid ;
wire merge1_split101_awready ;
wire [DWID-1:0] merge1_split101_wdata ;
wire [WSTRB-1:0] merge1_split101_wstrb ;
wire merge1_split101_wlast ;
wire merge1_split101_wvalid ;
wire merge1_split101_wready ;
wire [IDWID-1:0] merge1_split101_bid ;
wire [1:0] merge1_split101_bresp ;
wire merge1_split101_bvalid ;
wire merge1_split101_bready ;


wire [IDWID-1:0] split1_merge1_arid ;
wire [31:0] split1_merge1_araddr ;
wire [7:0] split1_merge1_arlen ;
wire [EXTRAS-1:0] split1_merge1_arextras ;
wire [1:0] split1_merge1_arburst ;
wire split1_merge1_arvalid ;
wire split1_merge1_arready ;
wire [IDWID-1:0] split1_merge1_rid ;
wire [DWID-1:0] split1_merge1_rdata ;
wire [1:0] split1_merge1_rresp ;
wire split1_merge1_rlast ;
wire split1_merge1_rvalid ;
wire split1_merge1_rready ;

wire [IDWID-1:0] split1_merge1_awid ;
wire [31:0] split1_merge1_awaddr ;
wire [7:0] split1_merge1_awlen ;
wire [EXTRAS-1:0] split1_merge1_awextras ;
wire [1:0] split1_merge1_awburst ;
wire split1_merge1_awvalid ;
wire split1_merge1_awready ;
wire [DWID-1:0] split1_merge1_wdata ;
wire [WSTRB-1:0] split1_merge1_wstrb ;
wire split1_merge1_wlast ;
wire split1_merge1_wvalid ;
wire split1_merge1_wready ;
wire [IDWID-1:0] split1_merge1_bid ;
wire [1:0] split1_merge1_bresp ;
wire split1_merge1_bvalid ;
wire split1_merge1_bready ;


wire [IDWID-1:0] split2_merge1_arid ;
wire [31:0] split2_merge1_araddr ;
wire [7:0] split2_merge1_arlen ;
wire [EXTRAS-1:0] split2_merge1_arextras ;
wire [1:0] split2_merge1_arburst ;
wire split2_merge1_arvalid ;
wire split2_merge1_arready ;
wire [IDWID-1:0] split2_merge1_rid ;
wire [DWID-1:0] split2_merge1_rdata ;
wire [1:0] split2_merge1_rresp ;
wire split2_merge1_rlast ;
wire split2_merge1_rvalid ;
wire split2_merge1_rready ;

wire [IDWID-1:0] split2_merge1_awid ;
wire [31:0] split2_merge1_awaddr ;
wire [7:0] split2_merge1_awlen ;
wire [EXTRAS-1:0] split2_merge1_awextras ;
wire [1:0] split2_merge1_awburst ;
wire split2_merge1_awvalid ;
wire split2_merge1_awready ;
wire [DWID-1:0] split2_merge1_wdata ;
wire [WSTRB-1:0] split2_merge1_wstrb ;
wire split2_merge1_wlast ;
wire split2_merge1_wvalid ;
wire split2_merge1_wready ;
wire [IDWID-1:0] split2_merge1_bid ;
wire [1:0] split2_merge1_bresp ;
wire split2_merge1_bvalid ;
wire split2_merge1_bready ;


wire [IDWID-1:0] split3_merge1_arid ;
wire [31:0] split3_merge1_araddr ;
wire [7:0] split3_merge1_arlen ;
wire [EXTRAS-1:0] split3_merge1_arextras ;
wire [1:0] split3_merge1_arburst ;
wire split3_merge1_arvalid ;
wire split3_merge1_arready ;
wire [IDWID-1:0] split3_merge1_rid ;
wire [DWID-1:0] split3_merge1_rdata ;
wire [1:0] split3_merge1_rresp ;
wire split3_merge1_rlast ;
wire split3_merge1_rvalid ;
wire split3_merge1_rready ;

wire [IDWID-1:0] split3_merge1_awid ;
wire [31:0] split3_merge1_awaddr ;
wire [7:0] split3_merge1_awlen ;
wire [EXTRAS-1:0] split3_merge1_awextras ;
wire [1:0] split3_merge1_awburst ;
wire split3_merge1_awvalid ;
wire split3_merge1_awready ;
wire [DWID-1:0] split3_merge1_wdata ;
wire [WSTRB-1:0] split3_merge1_wstrb ;
wire split3_merge1_wlast ;
wire split3_merge1_wvalid ;
wire split3_merge1_wready ;
wire [IDWID-1:0] split3_merge1_bid ;
wire [1:0] split3_merge1_bresp ;
wire split3_merge1_bvalid ;
wire split3_merge1_bready ;


axi_4_merger merge1 (
     .clk(clk),.rst_n(rst_n)
    ,.araddr(merge1_split101_araddr[31:0])
    ,.arburst(merge1_split101_arburst[1:0])
    ,.arextras(merge1_split101_arextras[(EXTRAS - 1):0])
    ,.arid(merge1_split101_arid[(IDWID - 1):0])
    ,.arlen(merge1_split101_arlen[7:0])
    ,.arready(merge1_split101_arready)
    ,.arvalid(merge1_split101_arvalid)
    ,.awaddr(merge1_split101_awaddr[31:0])
    ,.awburst(merge1_split101_awburst[1:0])
    ,.awextras(merge1_split101_awextras[(EXTRAS - 1):0])
    ,.awid(merge1_split101_awid[3:0])
    ,.awlen(merge1_split101_awlen[7:0])
    ,.awready(merge1_split101_awready)
    ,.awvalid(merge1_split101_awvalid)
    ,.bid(merge1_split101_bid[(IDWID - 1):0])
    ,.bready(merge1_split101_bready)
    ,.bresp(merge1_split101_bresp[1:0])
    ,.bvalid(merge1_split101_bvalid)
    ,.rid(merge1_split101_rid[(IDWID - 1):0])
    ,.rlast(merge1_split101_rlast)
    ,.rready(merge1_split101_rready)
    ,.rresp(merge1_split101_rresp[1:0])
    ,.rvalid(merge1_split101_rvalid)
    ,.rdata(merge1_split101_rdata[(DWID - 1):0])
    ,.wdata(merge1_split101_wdata[(DWID - 1):0])
    ,.wlast(merge1_split101_wlast)
    ,.wready(merge1_split101_wready)
    ,.wstrb(merge1_split101_wstrb[(WSTRB - 1):0])
    ,.wvalid(merge1_split101_wvalid)


    ,.a_araddr(split0_merge1_araddr[31:0])
    ,.a_arburst(split0_merge1_arburst[1:0])
    ,.a_arextras(split0_merge1_arextras[(EXTRAS - 1):0])
    ,.a_arid(split0_merge1_arid[(IDWID - 1):0])
    ,.a_arlen(split0_merge1_arlen[7:0])
    ,.a_arready(split0_merge1_arready)
    ,.a_arvalid(split0_merge1_arvalid)
    ,.a_awaddr(split0_merge1_awaddr[31:0])
    ,.a_awburst(split0_merge1_awburst[1:0])
    ,.a_awextras(split0_merge1_awextras[(EXTRAS - 1):0])
    ,.a_awid(split0_merge1_awid[(IDWID - 1):0])
    ,.a_awlen(split0_merge1_awlen[7:0])
    ,.a_awready(split0_merge1_awready)
    ,.a_awvalid(split0_merge1_awvalid)
    ,.a_bid(split0_merge1_bid[(IDWID - 1):0])
    ,.a_bready(split0_merge1_bready)
    ,.a_bresp(split0_merge1_bresp[1:0])
    ,.a_bvalid(split0_merge1_bvalid)
    ,.a_rdata(split0_merge1_rdata[(DWID - 1):0])
    ,.a_rid(split0_merge1_rid[(IDWID - 1):0])
    ,.a_rlast(split0_merge1_rlast)
    ,.a_rready(split0_merge1_rready)
    ,.a_rresp(split0_merge1_rresp[1:0])
    ,.a_rvalid(split0_merge1_rvalid)
    ,.a_wdata(split0_merge1_wdata[(DWID - 1):0])
    ,.a_wlast(split0_merge1_wlast)
    ,.a_wready(split0_merge1_wready)
    ,.a_wstrb(split0_merge1_wstrb[(WSTRB - 1):0])
    ,.a_wvalid(split0_merge1_wvalid)

    ,.b_araddr(split1_merge1_araddr[31:0])
    ,.b_arburst(split1_merge1_arburst[1:0])
    ,.b_arextras(split1_merge1_arextras[(EXTRAS - 1):0])
    ,.b_arid(split1_merge1_arid[(IDWID - 1):0])
    ,.b_arlen(split1_merge1_arlen[7:0])
    ,.b_arready(split1_merge1_arready)
    ,.b_arvalid(split1_merge1_arvalid)
    ,.b_awaddr(split1_merge1_awaddr[31:0])
    ,.b_awburst(split1_merge1_awburst[1:0])
    ,.b_awextras(split1_merge1_awextras[(EXTRAS - 1):0])
    ,.b_awid(split1_merge1_awid[(IDWID - 1):0])
    ,.b_awlen(split1_merge1_awlen[7:0])
    ,.b_awready(split1_merge1_awready)
    ,.b_awvalid(split1_merge1_awvalid)
    ,.b_bid(split1_merge1_bid[(IDWID - 1):0])
    ,.b_bready(split1_merge1_bready)
    ,.b_bresp(split1_merge1_bresp[1:0])
    ,.b_bvalid(split1_merge1_bvalid)
    ,.b_rdata(split1_merge1_rdata[(DWID - 1):0])
    ,.b_rid(split1_merge1_rid[(IDWID - 1):0])
    ,.b_rlast(split1_merge1_rlast)
    ,.b_rready(split1_merge1_rready)
    ,.b_rresp(split1_merge1_rresp[1:0])
    ,.b_rvalid(split1_merge1_rvalid)
    ,.b_wdata(split1_merge1_wdata[(DWID - 1):0])
    ,.b_wlast(split1_merge1_wlast)
    ,.b_wready(split1_merge1_wready)
    ,.b_wstrb(split1_merge1_wstrb[(WSTRB - 1):0])
    ,.b_wvalid(split1_merge1_wvalid)

    ,.c_araddr(split2_merge1_araddr[31:0])
    ,.c_arburst(split2_merge1_arburst[1:0])
    ,.c_arextras(split2_merge1_arextras[(EXTRAS - 1):0])
    ,.c_arid(split2_merge1_arid[(IDWID - 1):0])
    ,.c_arlen(split2_merge1_arlen[7:0])
    ,.c_arready(split2_merge1_arready)
    ,.c_arvalid(split2_merge1_arvalid)
    ,.c_awaddr(split2_merge1_awaddr[31:0])
    ,.c_awburst(split2_merge1_awburst[1:0])
    ,.c_awextras(split2_merge1_awextras[(EXTRAS - 1):0])
    ,.c_awid(split2_merge1_awid[(IDWID - 1):0])
    ,.c_awlen(split2_merge1_awlen[7:0])
    ,.c_awready(split2_merge1_awready)
    ,.c_awvalid(split2_merge1_awvalid)
    ,.c_bid(split2_merge1_bid[(IDWID - 1):0])
    ,.c_bready(split2_merge1_bready)
    ,.c_bresp(split2_merge1_bresp[1:0])
    ,.c_bvalid(split2_merge1_bvalid)
    ,.c_rdata(split2_merge1_rdata[(DWID - 1):0])
    ,.c_rid(split2_merge1_rid[(IDWID - 1):0])
    ,.c_rlast(split2_merge1_rlast)
    ,.c_rready(split2_merge1_rready)
    ,.c_rresp(split2_merge1_rresp[1:0])
    ,.c_rvalid(split2_merge1_rvalid)
    ,.c_wdata(split2_merge1_wdata[(DWID - 1):0])
    ,.c_wlast(split2_merge1_wlast)
    ,.c_wready(split2_merge1_wready)
    ,.c_wstrb(split2_merge1_wstrb[(WSTRB - 1):0])
    ,.c_wvalid(split2_merge1_wvalid)

    ,.d_araddr(split3_merge1_araddr[31:0])
    ,.d_arburst(split3_merge1_arburst[1:0])
    ,.d_arextras(split3_merge1_arextras[(EXTRAS - 1):0])
    ,.d_arid(split3_merge1_arid[(IDWID - 1):0])
    ,.d_arlen(split3_merge1_arlen[7:0])
    ,.d_arready(split3_merge1_arready)
    ,.d_arvalid(split3_merge1_arvalid)
    ,.d_awaddr(split3_merge1_awaddr[31:0])
    ,.d_awburst(split3_merge1_awburst[1:0])
    ,.d_awextras(split3_merge1_awextras[(EXTRAS - 1):0])
    ,.d_awid(split3_merge1_awid[(IDWID - 1):0])
    ,.d_awlen(split3_merge1_awlen[7:0])
    ,.d_awready(split3_merge1_awready)
    ,.d_awvalid(split3_merge1_awvalid)
    ,.d_bid(split3_merge1_bid[(IDWID - 1):0])
    ,.d_bready(split3_merge1_bready)
    ,.d_bresp(split3_merge1_bresp[1:0])
    ,.d_bvalid(split3_merge1_bvalid)
    ,.d_rdata(split3_merge1_rdata[(DWID - 1):0])
    ,.d_rid(split3_merge1_rid[(IDWID - 1):0])
    ,.d_rlast(split3_merge1_rlast)
    ,.d_rready(split3_merge1_rready)
    ,.d_rresp(split3_merge1_rresp[1:0])
    ,.d_rvalid(split3_merge1_rvalid)
    ,.d_wdata(split3_merge1_wdata[(DWID - 1):0])
    ,.d_wlast(split3_merge1_wlast)
    ,.d_wready(split3_merge1_wready)
    ,.d_wstrb(split3_merge1_wstrb[(WSTRB - 1):0])
    ,.d_wvalid(split3_merge1_wvalid)
);


wire [IDWID-1:0] merge2_split102_arid ;
wire [31:0] merge2_split102_araddr ;
wire [7:0] merge2_split102_arlen ;
wire [EXTRAS-1:0] merge2_split102_arextras ;
wire [1:0] merge2_split102_arburst ;
wire merge2_split102_arvalid ;
wire merge2_split102_arready ;
wire [IDWID-1:0] merge2_split102_rid ;
wire [DWID-1:0] merge2_split102_rdata ;
wire [1:0] merge2_split102_rresp ;
wire merge2_split102_rlast ;
wire merge2_split102_rvalid ;
wire merge2_split102_rready ;

wire [IDWID-1:0] merge2_split102_awid ;
wire [31:0] merge2_split102_awaddr ;
wire [7:0] merge2_split102_awlen ;
wire [EXTRAS-1:0] merge2_split102_awextras ;
wire [1:0] merge2_split102_awburst ;
wire merge2_split102_awvalid ;
wire merge2_split102_awready ;
wire [DWID-1:0] merge2_split102_wdata ;
wire [WSTRB-1:0] merge2_split102_wstrb ;
wire merge2_split102_wlast ;
wire merge2_split102_wvalid ;
wire merge2_split102_wready ;
wire [IDWID-1:0] merge2_split102_bid ;
wire [1:0] merge2_split102_bresp ;
wire merge2_split102_bvalid ;
wire merge2_split102_bready ;


wire [IDWID-1:0] split1_merge2_arid ;
wire [31:0] split1_merge2_araddr ;
wire [7:0] split1_merge2_arlen ;
wire [EXTRAS-1:0] split1_merge2_arextras ;
wire [1:0] split1_merge2_arburst ;
wire split1_merge2_arvalid ;
wire split1_merge2_arready ;
wire [IDWID-1:0] split1_merge2_rid ;
wire [DWID-1:0] split1_merge2_rdata ;
wire [1:0] split1_merge2_rresp ;
wire split1_merge2_rlast ;
wire split1_merge2_rvalid ;
wire split1_merge2_rready ;

wire [IDWID-1:0] split1_merge2_awid ;
wire [31:0] split1_merge2_awaddr ;
wire [7:0] split1_merge2_awlen ;
wire [EXTRAS-1:0] split1_merge2_awextras ;
wire [1:0] split1_merge2_awburst ;
wire split1_merge2_awvalid ;
wire split1_merge2_awready ;
wire [DWID-1:0] split1_merge2_wdata ;
wire [WSTRB-1:0] split1_merge2_wstrb ;
wire split1_merge2_wlast ;
wire split1_merge2_wvalid ;
wire split1_merge2_wready ;
wire [IDWID-1:0] split1_merge2_bid ;
wire [1:0] split1_merge2_bresp ;
wire split1_merge2_bvalid ;
wire split1_merge2_bready ;


wire [IDWID-1:0] split2_merge2_arid ;
wire [31:0] split2_merge2_araddr ;
wire [7:0] split2_merge2_arlen ;
wire [EXTRAS-1:0] split2_merge2_arextras ;
wire [1:0] split2_merge2_arburst ;
wire split2_merge2_arvalid ;
wire split2_merge2_arready ;
wire [IDWID-1:0] split2_merge2_rid ;
wire [DWID-1:0] split2_merge2_rdata ;
wire [1:0] split2_merge2_rresp ;
wire split2_merge2_rlast ;
wire split2_merge2_rvalid ;
wire split2_merge2_rready ;

wire [IDWID-1:0] split2_merge2_awid ;
wire [31:0] split2_merge2_awaddr ;
wire [7:0] split2_merge2_awlen ;
wire [EXTRAS-1:0] split2_merge2_awextras ;
wire [1:0] split2_merge2_awburst ;
wire split2_merge2_awvalid ;
wire split2_merge2_awready ;
wire [DWID-1:0] split2_merge2_wdata ;
wire [WSTRB-1:0] split2_merge2_wstrb ;
wire split2_merge2_wlast ;
wire split2_merge2_wvalid ;
wire split2_merge2_wready ;
wire [IDWID-1:0] split2_merge2_bid ;
wire [1:0] split2_merge2_bresp ;
wire split2_merge2_bvalid ;
wire split2_merge2_bready ;


wire [IDWID-1:0] split3_merge2_arid ;
wire [31:0] split3_merge2_araddr ;
wire [7:0] split3_merge2_arlen ;
wire [EXTRAS-1:0] split3_merge2_arextras ;
wire [1:0] split3_merge2_arburst ;
wire split3_merge2_arvalid ;
wire split3_merge2_arready ;
wire [IDWID-1:0] split3_merge2_rid ;
wire [DWID-1:0] split3_merge2_rdata ;
wire [1:0] split3_merge2_rresp ;
wire split3_merge2_rlast ;
wire split3_merge2_rvalid ;
wire split3_merge2_rready ;

wire [IDWID-1:0] split3_merge2_awid ;
wire [31:0] split3_merge2_awaddr ;
wire [7:0] split3_merge2_awlen ;
wire [EXTRAS-1:0] split3_merge2_awextras ;
wire [1:0] split3_merge2_awburst ;
wire split3_merge2_awvalid ;
wire split3_merge2_awready ;
wire [DWID-1:0] split3_merge2_wdata ;
wire [WSTRB-1:0] split3_merge2_wstrb ;
wire split3_merge2_wlast ;
wire split3_merge2_wvalid ;
wire split3_merge2_wready ;
wire [IDWID-1:0] split3_merge2_bid ;
wire [1:0] split3_merge2_bresp ;
wire split3_merge2_bvalid ;
wire split3_merge2_bready ;


axi_4_merger merge2 (
     .clk(clk),.rst_n(rst_n)
    ,.araddr(merge2_split102_araddr[31:0])
    ,.arburst(merge2_split102_arburst[1:0])
    ,.arextras(merge2_split102_arextras[(EXTRAS - 1):0])
    ,.arid(merge2_split102_arid[(IDWID - 1):0])
    ,.arlen(merge2_split102_arlen[7:0])
    ,.arready(merge2_split102_arready)
    ,.arvalid(merge2_split102_arvalid)
    ,.awaddr(merge2_split102_awaddr[31:0])
    ,.awburst(merge2_split102_awburst[1:0])
    ,.awextras(merge2_split102_awextras[(EXTRAS - 1):0])
    ,.awid(merge2_split102_awid[3:0])
    ,.awlen(merge2_split102_awlen[7:0])
    ,.awready(merge2_split102_awready)
    ,.awvalid(merge2_split102_awvalid)
    ,.bid(merge2_split102_bid[(IDWID - 1):0])
    ,.bready(merge2_split102_bready)
    ,.bresp(merge2_split102_bresp[1:0])
    ,.bvalid(merge2_split102_bvalid)
    ,.rid(merge2_split102_rid[(IDWID - 1):0])
    ,.rlast(merge2_split102_rlast)
    ,.rready(merge2_split102_rready)
    ,.rresp(merge2_split102_rresp[1:0])
    ,.rvalid(merge2_split102_rvalid)
    ,.rdata(merge2_split102_rdata[(DWID - 1):0])
    ,.wdata(merge2_split102_wdata[(DWID - 1):0])
    ,.wlast(merge2_split102_wlast)
    ,.wready(merge2_split102_wready)
    ,.wstrb(merge2_split102_wstrb[(WSTRB - 1):0])
    ,.wvalid(merge2_split102_wvalid)


    ,.a_araddr(split0_merge2_araddr[31:0])
    ,.a_arburst(split0_merge2_arburst[1:0])
    ,.a_arextras(split0_merge2_arextras[(EXTRAS - 1):0])
    ,.a_arid(split0_merge2_arid[(IDWID - 1):0])
    ,.a_arlen(split0_merge2_arlen[7:0])
    ,.a_arready(split0_merge2_arready)
    ,.a_arvalid(split0_merge2_arvalid)
    ,.a_awaddr(split0_merge2_awaddr[31:0])
    ,.a_awburst(split0_merge2_awburst[1:0])
    ,.a_awextras(split0_merge2_awextras[(EXTRAS - 1):0])
    ,.a_awid(split0_merge2_awid[(IDWID - 1):0])
    ,.a_awlen(split0_merge2_awlen[7:0])
    ,.a_awready(split0_merge2_awready)
    ,.a_awvalid(split0_merge2_awvalid)
    ,.a_bid(split0_merge2_bid[(IDWID - 1):0])
    ,.a_bready(split0_merge2_bready)
    ,.a_bresp(split0_merge2_bresp[1:0])
    ,.a_bvalid(split0_merge2_bvalid)
    ,.a_rdata(split0_merge2_rdata[(DWID - 1):0])
    ,.a_rid(split0_merge2_rid[(IDWID - 1):0])
    ,.a_rlast(split0_merge2_rlast)
    ,.a_rready(split0_merge2_rready)
    ,.a_rresp(split0_merge2_rresp[1:0])
    ,.a_rvalid(split0_merge2_rvalid)
    ,.a_wdata(split0_merge2_wdata[(DWID - 1):0])
    ,.a_wlast(split0_merge2_wlast)
    ,.a_wready(split0_merge2_wready)
    ,.a_wstrb(split0_merge2_wstrb[(WSTRB - 1):0])
    ,.a_wvalid(split0_merge2_wvalid)

    ,.b_araddr(split1_merge2_araddr[31:0])
    ,.b_arburst(split1_merge2_arburst[1:0])
    ,.b_arextras(split1_merge2_arextras[(EXTRAS - 1):0])
    ,.b_arid(split1_merge2_arid[(IDWID - 1):0])
    ,.b_arlen(split1_merge2_arlen[7:0])
    ,.b_arready(split1_merge2_arready)
    ,.b_arvalid(split1_merge2_arvalid)
    ,.b_awaddr(split1_merge2_awaddr[31:0])
    ,.b_awburst(split1_merge2_awburst[1:0])
    ,.b_awextras(split1_merge2_awextras[(EXTRAS - 1):0])
    ,.b_awid(split1_merge2_awid[(IDWID - 1):0])
    ,.b_awlen(split1_merge2_awlen[7:0])
    ,.b_awready(split1_merge2_awready)
    ,.b_awvalid(split1_merge2_awvalid)
    ,.b_bid(split1_merge2_bid[(IDWID - 1):0])
    ,.b_bready(split1_merge2_bready)
    ,.b_bresp(split1_merge2_bresp[1:0])
    ,.b_bvalid(split1_merge2_bvalid)
    ,.b_rdata(split1_merge2_rdata[(DWID - 1):0])
    ,.b_rid(split1_merge2_rid[(IDWID - 1):0])
    ,.b_rlast(split1_merge2_rlast)
    ,.b_rready(split1_merge2_rready)
    ,.b_rresp(split1_merge2_rresp[1:0])
    ,.b_rvalid(split1_merge2_rvalid)
    ,.b_wdata(split1_merge2_wdata[(DWID - 1):0])
    ,.b_wlast(split1_merge2_wlast)
    ,.b_wready(split1_merge2_wready)
    ,.b_wstrb(split1_merge2_wstrb[(WSTRB - 1):0])
    ,.b_wvalid(split1_merge2_wvalid)

    ,.c_araddr(split2_merge2_araddr[31:0])
    ,.c_arburst(split2_merge2_arburst[1:0])
    ,.c_arextras(split2_merge2_arextras[(EXTRAS - 1):0])
    ,.c_arid(split2_merge2_arid[(IDWID - 1):0])
    ,.c_arlen(split2_merge2_arlen[7:0])
    ,.c_arready(split2_merge2_arready)
    ,.c_arvalid(split2_merge2_arvalid)
    ,.c_awaddr(split2_merge2_awaddr[31:0])
    ,.c_awburst(split2_merge2_awburst[1:0])
    ,.c_awextras(split2_merge2_awextras[(EXTRAS - 1):0])
    ,.c_awid(split2_merge2_awid[(IDWID - 1):0])
    ,.c_awlen(split2_merge2_awlen[7:0])
    ,.c_awready(split2_merge2_awready)
    ,.c_awvalid(split2_merge2_awvalid)
    ,.c_bid(split2_merge2_bid[(IDWID - 1):0])
    ,.c_bready(split2_merge2_bready)
    ,.c_bresp(split2_merge2_bresp[1:0])
    ,.c_bvalid(split2_merge2_bvalid)
    ,.c_rdata(split2_merge2_rdata[(DWID - 1):0])
    ,.c_rid(split2_merge2_rid[(IDWID - 1):0])
    ,.c_rlast(split2_merge2_rlast)
    ,.c_rready(split2_merge2_rready)
    ,.c_rresp(split2_merge2_rresp[1:0])
    ,.c_rvalid(split2_merge2_rvalid)
    ,.c_wdata(split2_merge2_wdata[(DWID - 1):0])
    ,.c_wlast(split2_merge2_wlast)
    ,.c_wready(split2_merge2_wready)
    ,.c_wstrb(split2_merge2_wstrb[(WSTRB - 1):0])
    ,.c_wvalid(split2_merge2_wvalid)

    ,.d_araddr(split3_merge2_araddr[31:0])
    ,.d_arburst(split3_merge2_arburst[1:0])
    ,.d_arextras(split3_merge2_arextras[(EXTRAS - 1):0])
    ,.d_arid(split3_merge2_arid[(IDWID - 1):0])
    ,.d_arlen(split3_merge2_arlen[7:0])
    ,.d_arready(split3_merge2_arready)
    ,.d_arvalid(split3_merge2_arvalid)
    ,.d_awaddr(split3_merge2_awaddr[31:0])
    ,.d_awburst(split3_merge2_awburst[1:0])
    ,.d_awextras(split3_merge2_awextras[(EXTRAS - 1):0])
    ,.d_awid(split3_merge2_awid[(IDWID - 1):0])
    ,.d_awlen(split3_merge2_awlen[7:0])
    ,.d_awready(split3_merge2_awready)
    ,.d_awvalid(split3_merge2_awvalid)
    ,.d_bid(split3_merge2_bid[(IDWID - 1):0])
    ,.d_bready(split3_merge2_bready)
    ,.d_bresp(split3_merge2_bresp[1:0])
    ,.d_bvalid(split3_merge2_bvalid)
    ,.d_rdata(split3_merge2_rdata[(DWID - 1):0])
    ,.d_rid(split3_merge2_rid[(IDWID - 1):0])
    ,.d_rlast(split3_merge2_rlast)
    ,.d_rready(split3_merge2_rready)
    ,.d_rresp(split3_merge2_rresp[1:0])
    ,.d_rvalid(split3_merge2_rvalid)
    ,.d_wdata(split3_merge2_wdata[(DWID - 1):0])
    ,.d_wlast(split3_merge2_wlast)
    ,.d_wready(split3_merge2_wready)
    ,.d_wstrb(split3_merge2_wstrb[(WSTRB - 1):0])
    ,.d_wvalid(split3_merge2_wvalid)
);


wire [IDWID-1:0] merge3_split103_arid ;
wire [31:0] merge3_split103_araddr ;
wire [7:0] merge3_split103_arlen ;
wire [EXTRAS-1:0] merge3_split103_arextras ;
wire [1:0] merge3_split103_arburst ;
wire merge3_split103_arvalid ;
wire merge3_split103_arready ;
wire [IDWID-1:0] merge3_split103_rid ;
wire [DWID-1:0] merge3_split103_rdata ;
wire [1:0] merge3_split103_rresp ;
wire merge3_split103_rlast ;
wire merge3_split103_rvalid ;
wire merge3_split103_rready ;

wire [IDWID-1:0] merge3_split103_awid ;
wire [31:0] merge3_split103_awaddr ;
wire [7:0] merge3_split103_awlen ;
wire [EXTRAS-1:0] merge3_split103_awextras ;
wire [1:0] merge3_split103_awburst ;
wire merge3_split103_awvalid ;
wire merge3_split103_awready ;
wire [DWID-1:0] merge3_split103_wdata ;
wire [WSTRB-1:0] merge3_split103_wstrb ;
wire merge3_split103_wlast ;
wire merge3_split103_wvalid ;
wire merge3_split103_wready ;
wire [IDWID-1:0] merge3_split103_bid ;
wire [1:0] merge3_split103_bresp ;
wire merge3_split103_bvalid ;
wire merge3_split103_bready ;


wire [IDWID-1:0] split1_merge3_arid ;
wire [31:0] split1_merge3_araddr ;
wire [7:0] split1_merge3_arlen ;
wire [EXTRAS-1:0] split1_merge3_arextras ;
wire [1:0] split1_merge3_arburst ;
wire split1_merge3_arvalid ;
wire split1_merge3_arready ;
wire [IDWID-1:0] split1_merge3_rid ;
wire [DWID-1:0] split1_merge3_rdata ;
wire [1:0] split1_merge3_rresp ;
wire split1_merge3_rlast ;
wire split1_merge3_rvalid ;
wire split1_merge3_rready ;

wire [IDWID-1:0] split1_merge3_awid ;
wire [31:0] split1_merge3_awaddr ;
wire [7:0] split1_merge3_awlen ;
wire [EXTRAS-1:0] split1_merge3_awextras ;
wire [1:0] split1_merge3_awburst ;
wire split1_merge3_awvalid ;
wire split1_merge3_awready ;
wire [DWID-1:0] split1_merge3_wdata ;
wire [WSTRB-1:0] split1_merge3_wstrb ;
wire split1_merge3_wlast ;
wire split1_merge3_wvalid ;
wire split1_merge3_wready ;
wire [IDWID-1:0] split1_merge3_bid ;
wire [1:0] split1_merge3_bresp ;
wire split1_merge3_bvalid ;
wire split1_merge3_bready ;


wire [IDWID-1:0] split2_merge3_arid ;
wire [31:0] split2_merge3_araddr ;
wire [7:0] split2_merge3_arlen ;
wire [EXTRAS-1:0] split2_merge3_arextras ;
wire [1:0] split2_merge3_arburst ;
wire split2_merge3_arvalid ;
wire split2_merge3_arready ;
wire [IDWID-1:0] split2_merge3_rid ;
wire [DWID-1:0] split2_merge3_rdata ;
wire [1:0] split2_merge3_rresp ;
wire split2_merge3_rlast ;
wire split2_merge3_rvalid ;
wire split2_merge3_rready ;

wire [IDWID-1:0] split2_merge3_awid ;
wire [31:0] split2_merge3_awaddr ;
wire [7:0] split2_merge3_awlen ;
wire [EXTRAS-1:0] split2_merge3_awextras ;
wire [1:0] split2_merge3_awburst ;
wire split2_merge3_awvalid ;
wire split2_merge3_awready ;
wire [DWID-1:0] split2_merge3_wdata ;
wire [WSTRB-1:0] split2_merge3_wstrb ;
wire split2_merge3_wlast ;
wire split2_merge3_wvalid ;
wire split2_merge3_wready ;
wire [IDWID-1:0] split2_merge3_bid ;
wire [1:0] split2_merge3_bresp ;
wire split2_merge3_bvalid ;
wire split2_merge3_bready ;


wire [IDWID-1:0] split3_merge3_arid ;
wire [31:0] split3_merge3_araddr ;
wire [7:0] split3_merge3_arlen ;
wire [EXTRAS-1:0] split3_merge3_arextras ;
wire [1:0] split3_merge3_arburst ;
wire split3_merge3_arvalid ;
wire split3_merge3_arready ;
wire [IDWID-1:0] split3_merge3_rid ;
wire [DWID-1:0] split3_merge3_rdata ;
wire [1:0] split3_merge3_rresp ;
wire split3_merge3_rlast ;
wire split3_merge3_rvalid ;
wire split3_merge3_rready ;

wire [IDWID-1:0] split3_merge3_awid ;
wire [31:0] split3_merge3_awaddr ;
wire [7:0] split3_merge3_awlen ;
wire [EXTRAS-1:0] split3_merge3_awextras ;
wire [1:0] split3_merge3_awburst ;
wire split3_merge3_awvalid ;
wire split3_merge3_awready ;
wire [DWID-1:0] split3_merge3_wdata ;
wire [WSTRB-1:0] split3_merge3_wstrb ;
wire split3_merge3_wlast ;
wire split3_merge3_wvalid ;
wire split3_merge3_wready ;
wire [IDWID-1:0] split3_merge3_bid ;
wire [1:0] split3_merge3_bresp ;
wire split3_merge3_bvalid ;
wire split3_merge3_bready ;


axi_4_merger merge3 (
     .clk(clk),.rst_n(rst_n)
    ,.araddr(merge3_split103_araddr[31:0])
    ,.arburst(merge3_split103_arburst[1:0])
    ,.arextras(merge3_split103_arextras[(EXTRAS - 1):0])
    ,.arid(merge3_split103_arid[(IDWID - 1):0])
    ,.arlen(merge3_split103_arlen[7:0])
    ,.arready(merge3_split103_arready)
    ,.arvalid(merge3_split103_arvalid)
    ,.awaddr(merge3_split103_awaddr[31:0])
    ,.awburst(merge3_split103_awburst[1:0])
    ,.awextras(merge3_split103_awextras[(EXTRAS - 1):0])
    ,.awid(merge3_split103_awid[3:0])
    ,.awlen(merge3_split103_awlen[7:0])
    ,.awready(merge3_split103_awready)
    ,.awvalid(merge3_split103_awvalid)
    ,.bid(merge3_split103_bid[(IDWID - 1):0])
    ,.bready(merge3_split103_bready)
    ,.bresp(merge3_split103_bresp[1:0])
    ,.bvalid(merge3_split103_bvalid)
    ,.rid(merge3_split103_rid[(IDWID - 1):0])
    ,.rlast(merge3_split103_rlast)
    ,.rready(merge3_split103_rready)
    ,.rresp(merge3_split103_rresp[1:0])
    ,.rvalid(merge3_split103_rvalid)
    ,.rdata(merge3_split103_rdata[(DWID - 1):0])
    ,.wdata(merge3_split103_wdata[(DWID - 1):0])
    ,.wlast(merge3_split103_wlast)
    ,.wready(merge3_split103_wready)
    ,.wstrb(merge3_split103_wstrb[(WSTRB - 1):0])
    ,.wvalid(merge3_split103_wvalid)


    ,.a_araddr(split0_merge3_araddr[31:0])
    ,.a_arburst(split0_merge3_arburst[1:0])
    ,.a_arextras(split0_merge3_arextras[(EXTRAS - 1):0])
    ,.a_arid(split0_merge3_arid[(IDWID - 1):0])
    ,.a_arlen(split0_merge3_arlen[7:0])
    ,.a_arready(split0_merge3_arready)
    ,.a_arvalid(split0_merge3_arvalid)
    ,.a_awaddr(split0_merge3_awaddr[31:0])
    ,.a_awburst(split0_merge3_awburst[1:0])
    ,.a_awextras(split0_merge3_awextras[(EXTRAS - 1):0])
    ,.a_awid(split0_merge3_awid[(IDWID - 1):0])
    ,.a_awlen(split0_merge3_awlen[7:0])
    ,.a_awready(split0_merge3_awready)
    ,.a_awvalid(split0_merge3_awvalid)
    ,.a_bid(split0_merge3_bid[(IDWID - 1):0])
    ,.a_bready(split0_merge3_bready)
    ,.a_bresp(split0_merge3_bresp[1:0])
    ,.a_bvalid(split0_merge3_bvalid)
    ,.a_rdata(split0_merge3_rdata[(DWID - 1):0])
    ,.a_rid(split0_merge3_rid[(IDWID - 1):0])
    ,.a_rlast(split0_merge3_rlast)
    ,.a_rready(split0_merge3_rready)
    ,.a_rresp(split0_merge3_rresp[1:0])
    ,.a_rvalid(split0_merge3_rvalid)
    ,.a_wdata(split0_merge3_wdata[(DWID - 1):0])
    ,.a_wlast(split0_merge3_wlast)
    ,.a_wready(split0_merge3_wready)
    ,.a_wstrb(split0_merge3_wstrb[(WSTRB - 1):0])
    ,.a_wvalid(split0_merge3_wvalid)

    ,.b_araddr(split1_merge3_araddr[31:0])
    ,.b_arburst(split1_merge3_arburst[1:0])
    ,.b_arextras(split1_merge3_arextras[(EXTRAS - 1):0])
    ,.b_arid(split1_merge3_arid[(IDWID - 1):0])
    ,.b_arlen(split1_merge3_arlen[7:0])
    ,.b_arready(split1_merge3_arready)
    ,.b_arvalid(split1_merge3_arvalid)
    ,.b_awaddr(split1_merge3_awaddr[31:0])
    ,.b_awburst(split1_merge3_awburst[1:0])
    ,.b_awextras(split1_merge3_awextras[(EXTRAS - 1):0])
    ,.b_awid(split1_merge3_awid[(IDWID - 1):0])
    ,.b_awlen(split1_merge3_awlen[7:0])
    ,.b_awready(split1_merge3_awready)
    ,.b_awvalid(split1_merge3_awvalid)
    ,.b_bid(split1_merge3_bid[(IDWID - 1):0])
    ,.b_bready(split1_merge3_bready)
    ,.b_bresp(split1_merge3_bresp[1:0])
    ,.b_bvalid(split1_merge3_bvalid)
    ,.b_rdata(split1_merge3_rdata[(DWID - 1):0])
    ,.b_rid(split1_merge3_rid[(IDWID - 1):0])
    ,.b_rlast(split1_merge3_rlast)
    ,.b_rready(split1_merge3_rready)
    ,.b_rresp(split1_merge3_rresp[1:0])
    ,.b_rvalid(split1_merge3_rvalid)
    ,.b_wdata(split1_merge3_wdata[(DWID - 1):0])
    ,.b_wlast(split1_merge3_wlast)
    ,.b_wready(split1_merge3_wready)
    ,.b_wstrb(split1_merge3_wstrb[(WSTRB - 1):0])
    ,.b_wvalid(split1_merge3_wvalid)

    ,.c_araddr(split2_merge3_araddr[31:0])
    ,.c_arburst(split2_merge3_arburst[1:0])
    ,.c_arextras(split2_merge3_arextras[(EXTRAS - 1):0])
    ,.c_arid(split2_merge3_arid[(IDWID - 1):0])
    ,.c_arlen(split2_merge3_arlen[7:0])
    ,.c_arready(split2_merge3_arready)
    ,.c_arvalid(split2_merge3_arvalid)
    ,.c_awaddr(split2_merge3_awaddr[31:0])
    ,.c_awburst(split2_merge3_awburst[1:0])
    ,.c_awextras(split2_merge3_awextras[(EXTRAS - 1):0])
    ,.c_awid(split2_merge3_awid[(IDWID - 1):0])
    ,.c_awlen(split2_merge3_awlen[7:0])
    ,.c_awready(split2_merge3_awready)
    ,.c_awvalid(split2_merge3_awvalid)
    ,.c_bid(split2_merge3_bid[(IDWID - 1):0])
    ,.c_bready(split2_merge3_bready)
    ,.c_bresp(split2_merge3_bresp[1:0])
    ,.c_bvalid(split2_merge3_bvalid)
    ,.c_rdata(split2_merge3_rdata[(DWID - 1):0])
    ,.c_rid(split2_merge3_rid[(IDWID - 1):0])
    ,.c_rlast(split2_merge3_rlast)
    ,.c_rready(split2_merge3_rready)
    ,.c_rresp(split2_merge3_rresp[1:0])
    ,.c_rvalid(split2_merge3_rvalid)
    ,.c_wdata(split2_merge3_wdata[(DWID - 1):0])
    ,.c_wlast(split2_merge3_wlast)
    ,.c_wready(split2_merge3_wready)
    ,.c_wstrb(split2_merge3_wstrb[(WSTRB - 1):0])
    ,.c_wvalid(split2_merge3_wvalid)

    ,.d_araddr(split3_merge3_araddr[31:0])
    ,.d_arburst(split3_merge3_arburst[1:0])
    ,.d_arextras(split3_merge3_arextras[(EXTRAS - 1):0])
    ,.d_arid(split3_merge3_arid[(IDWID - 1):0])
    ,.d_arlen(split3_merge3_arlen[7:0])
    ,.d_arready(split3_merge3_arready)
    ,.d_arvalid(split3_merge3_arvalid)
    ,.d_awaddr(split3_merge3_awaddr[31:0])
    ,.d_awburst(split3_merge3_awburst[1:0])
    ,.d_awextras(split3_merge3_awextras[(EXTRAS - 1):0])
    ,.d_awid(split3_merge3_awid[(IDWID - 1):0])
    ,.d_awlen(split3_merge3_awlen[7:0])
    ,.d_awready(split3_merge3_awready)
    ,.d_awvalid(split3_merge3_awvalid)
    ,.d_bid(split3_merge3_bid[(IDWID - 1):0])
    ,.d_bready(split3_merge3_bready)
    ,.d_bresp(split3_merge3_bresp[1:0])
    ,.d_bvalid(split3_merge3_bvalid)
    ,.d_rdata(split3_merge3_rdata[(DWID - 1):0])
    ,.d_rid(split3_merge3_rid[(IDWID - 1):0])
    ,.d_rlast(split3_merge3_rlast)
    ,.d_rready(split3_merge3_rready)
    ,.d_rresp(split3_merge3_rresp[1:0])
    ,.d_rvalid(split3_merge3_rvalid)
    ,.d_wdata(split3_merge3_wdata[(DWID - 1):0])
    ,.d_wlast(split3_merge3_wlast)
    ,.d_wready(split3_merge3_wready)
    ,.d_wstrb(split3_merge3_wstrb[(WSTRB - 1):0])
    ,.d_wvalid(split3_merge3_wvalid)
);


axi_4_splitter split1 (
     .clk(clk) ,.rst_n(rst_n)

    ,.araddr(mst1_araddr[31:0])
    ,.arburst(mst1_arburst[1:0])
    ,.arextras(mst1_arextras[(EXTRAS - 1):0])
    ,.arid(mst1_arid[(IDWID - 1):0])
    ,.arlen(mst1_arlen[7:0])
    ,.arready(mst1_arready)
    ,.arvalid(mst1_arvalid)
    ,.awaddr(mst1_awaddr[31:0])
    ,.awburst(mst1_awburst[1:0])
    ,.awextras(mst1_awextras[(EXTRAS - 1):0])
    ,.awid(mst1_awid[3:0])
    ,.awlen(mst1_awlen[7:0])
    ,.awready(mst1_awready)
    ,.awvalid(mst1_awvalid)
    ,.bid(mst1_bid[(IDWID - 1):0])
    ,.bready(mst1_bready)
    ,.bresp(mst1_bresp[1:0])
    ,.bvalid(mst1_bvalid)
    ,.rdata(mst1_rdata[(DWID - 1):0])
    ,.rid(mst1_rid[(IDWID - 1):0])
    ,.rlast(mst1_rlast)
    ,.rready(mst1_rready)
    ,.rresp(mst1_rresp[1:0])
    ,.rvalid(mst1_rvalid)
    ,.wdata(mst1_wdata[(DWID - 1):0])
    ,.wlast(mst1_wlast)
    ,.wready(mst1_wready)
    ,.wstrb(mst1_wstrb[(WSTRB - 1):0])
    ,.wvalid(mst1_wvalid)

    ,.a_araddr(split1_merge0_araddr[31:0])
    ,.a_arburst(split1_merge0_arburst[1:0])
    ,.a_arextras(split1_merge0_arextras[(EXTRAS - 1):0])
    ,.a_arid(split1_merge0_arid[(IDWID - 1):0])
    ,.a_arlen(split1_merge0_arlen[7:0])
    ,.a_arready(split1_merge0_arready)
    ,.a_arvalid(split1_merge0_arvalid)
    ,.a_awaddr(split1_merge0_awaddr[31:0])
    ,.a_awburst(split1_merge0_awburst[1:0])
    ,.a_awextras(split1_merge0_awextras[(EXTRAS - 1):0])
    ,.a_awid(split1_merge0_awid[(IDWID - 1):0])
    ,.a_awlen(split1_merge0_awlen[7:0])
    ,.a_awready(split1_merge0_awready)
    ,.a_awvalid(split1_merge0_awvalid)
    ,.a_bid(split1_merge0_bid[(IDWID - 1):0])
    ,.a_bready(split1_merge0_bready)
    ,.a_bresp(split1_merge0_bresp[1:0])
    ,.a_bvalid(split1_merge0_bvalid)
    ,.a_rdata(split1_merge0_rdata[(DWID - 1):0])
    ,.a_rid(split1_merge0_rid[(IDWID - 1):0])
    ,.a_rlast(split1_merge0_rlast)
    ,.a_rready(split1_merge0_rready)
    ,.a_rresp(split1_merge0_rresp[1:0])
    ,.a_rvalid(split1_merge0_rvalid)
    ,.a_wdata(split1_merge0_wdata[(DWID - 1):0])
    ,.a_wlast(split1_merge0_wlast)
    ,.a_wready(split1_merge0_wready)
    ,.a_wstrb(split1_merge0_wstrb[(WSTRB - 1):0])
    ,.a_wvalid(split1_merge0_wvalid)
    ,.b_araddr(split1_merge1_araddr[31:0])
    ,.b_arburst(split1_merge1_arburst[1:0])
    ,.b_arextras(split1_merge1_arextras[(EXTRAS - 1):0])
    ,.b_arid(split1_merge1_arid[(IDWID - 1):0])
    ,.b_arlen(split1_merge1_arlen[7:0])
    ,.b_arready(split1_merge1_arready)
    ,.b_arvalid(split1_merge1_arvalid)
    ,.b_awaddr(split1_merge1_awaddr[31:0])
    ,.b_awburst(split1_merge1_awburst[1:0])
    ,.b_awextras(split1_merge1_awextras[(EXTRAS - 1):0])
    ,.b_awid(split1_merge1_awid[(IDWID - 1):0])
    ,.b_awlen(split1_merge1_awlen[7:0])
    ,.b_awready(split1_merge1_awready)
    ,.b_awvalid(split1_merge1_awvalid)
    ,.b_bid(split1_merge1_bid[(IDWID - 1):0])
    ,.b_bready(split1_merge1_bready)
    ,.b_bresp(split1_merge1_bresp[1:0])
    ,.b_bvalid(split1_merge1_bvalid)
    ,.b_rdata(split1_merge1_rdata[(DWID - 1):0])
    ,.b_rid(split1_merge1_rid[(IDWID - 1):0])
    ,.b_rlast(split1_merge1_rlast)
    ,.b_rready(split1_merge1_rready)
    ,.b_rresp(split1_merge1_rresp[1:0])
    ,.b_rvalid(split1_merge1_rvalid)
    ,.b_wdata(split1_merge1_wdata[(DWID - 1):0])
    ,.b_wlast(split1_merge1_wlast)
    ,.b_wready(split1_merge1_wready)
    ,.b_wstrb(split1_merge1_wstrb[(WSTRB - 1):0])
    ,.b_wvalid(split1_merge1_wvalid)
    ,.c_araddr(split1_merge2_araddr[31:0])
    ,.c_arburst(split1_merge2_arburst[1:0])
    ,.c_arextras(split1_merge2_arextras[(EXTRAS - 1):0])
    ,.c_arid(split1_merge2_arid[(IDWID - 1):0])
    ,.c_arlen(split1_merge2_arlen[7:0])
    ,.c_arready(split1_merge2_arready)
    ,.c_arvalid(split1_merge2_arvalid)
    ,.c_awaddr(split1_merge2_awaddr[31:0])
    ,.c_awburst(split1_merge2_awburst[1:0])
    ,.c_awextras(split1_merge2_awextras[(EXTRAS - 1):0])
    ,.c_awid(split1_merge2_awid[(IDWID - 1):0])
    ,.c_awlen(split1_merge2_awlen[7:0])
    ,.c_awready(split1_merge2_awready)
    ,.c_awvalid(split1_merge2_awvalid)
    ,.c_bid(split1_merge2_bid[(IDWID - 1):0])
    ,.c_bready(split1_merge2_bready)
    ,.c_bresp(split1_merge2_bresp[1:0])
    ,.c_bvalid(split1_merge2_bvalid)
    ,.c_rdata(split1_merge2_rdata[(DWID - 1):0])
    ,.c_rid(split1_merge2_rid[(IDWID - 1):0])
    ,.c_rlast(split1_merge2_rlast)
    ,.c_rready(split1_merge2_rready)
    ,.c_rresp(split1_merge2_rresp[1:0])
    ,.c_rvalid(split1_merge2_rvalid)
    ,.c_wdata(split1_merge2_wdata[(DWID - 1):0])
    ,.c_wlast(split1_merge2_wlast)
    ,.c_wready(split1_merge2_wready)
    ,.c_wstrb(split1_merge2_wstrb[(WSTRB - 1):0])
    ,.c_wvalid(split1_merge2_wvalid)
    ,.d_araddr(split1_merge3_araddr[31:0])
    ,.d_arburst(split1_merge3_arburst[1:0])
    ,.d_arextras(split1_merge3_arextras[(EXTRAS - 1):0])
    ,.d_arid(split1_merge3_arid[(IDWID - 1):0])
    ,.d_arlen(split1_merge3_arlen[7:0])
    ,.d_arready(split1_merge3_arready)
    ,.d_arvalid(split1_merge3_arvalid)
    ,.d_awaddr(split1_merge3_awaddr[31:0])
    ,.d_awburst(split1_merge3_awburst[1:0])
    ,.d_awextras(split1_merge3_awextras[(EXTRAS - 1):0])
    ,.d_awid(split1_merge3_awid[(IDWID - 1):0])
    ,.d_awlen(split1_merge3_awlen[7:0])
    ,.d_awready(split1_merge3_awready)
    ,.d_awvalid(split1_merge3_awvalid)
    ,.d_bid(split1_merge3_bid[(IDWID - 1):0])
    ,.d_bready(split1_merge3_bready)
    ,.d_bresp(split1_merge3_bresp[1:0])
    ,.d_bvalid(split1_merge3_bvalid)
    ,.d_rdata(split1_merge3_rdata[(DWID - 1):0])
    ,.d_rid(split1_merge3_rid[(IDWID - 1):0])
    ,.d_rlast(split1_merge3_rlast)
    ,.d_rready(split1_merge3_rready)
    ,.d_rresp(split1_merge3_rresp[1:0])
    ,.d_rvalid(split1_merge3_rvalid)
    ,.d_wdata(split1_merge3_wdata[(DWID - 1):0])
    ,.d_wlast(split1_merge3_wlast)
    ,.d_wready(split1_merge3_wready)
    ,.d_wstrb(split1_merge3_wstrb[(WSTRB - 1):0])
    ,.d_wvalid(split1_merge3_wvalid)

);

axi_4_splitter split2 (
     .clk(clk) ,.rst_n(rst_n)

    ,.araddr(mst2_araddr[31:0])
    ,.arburst(mst2_arburst[1:0])
    ,.arextras(mst2_arextras[(EXTRAS - 1):0])
    ,.arid(mst2_arid[(IDWID - 1):0])
    ,.arlen(mst2_arlen[7:0])
    ,.arready(mst2_arready)
    ,.arvalid(mst2_arvalid)
    ,.awaddr(mst2_awaddr[31:0])
    ,.awburst(mst2_awburst[1:0])
    ,.awextras(mst2_awextras[(EXTRAS - 1):0])
    ,.awid(mst2_awid[3:0])
    ,.awlen(mst2_awlen[7:0])
    ,.awready(mst2_awready)
    ,.awvalid(mst2_awvalid)
    ,.bid(mst2_bid[(IDWID - 1):0])
    ,.bready(mst2_bready)
    ,.bresp(mst2_bresp[1:0])
    ,.bvalid(mst2_bvalid)
    ,.rdata(mst2_rdata[(DWID - 1):0])
    ,.rid(mst2_rid[(IDWID - 1):0])
    ,.rlast(mst2_rlast)
    ,.rready(mst2_rready)
    ,.rresp(mst2_rresp[1:0])
    ,.rvalid(mst2_rvalid)
    ,.wdata(mst2_wdata[(DWID - 1):0])
    ,.wlast(mst2_wlast)
    ,.wready(mst2_wready)
    ,.wstrb(mst2_wstrb[(WSTRB - 1):0])
    ,.wvalid(mst2_wvalid)

    ,.a_araddr(split2_merge0_araddr[31:0])
    ,.a_arburst(split2_merge0_arburst[1:0])
    ,.a_arextras(split2_merge0_arextras[(EXTRAS - 1):0])
    ,.a_arid(split2_merge0_arid[(IDWID - 1):0])
    ,.a_arlen(split2_merge0_arlen[7:0])
    ,.a_arready(split2_merge0_arready)
    ,.a_arvalid(split2_merge0_arvalid)
    ,.a_awaddr(split2_merge0_awaddr[31:0])
    ,.a_awburst(split2_merge0_awburst[1:0])
    ,.a_awextras(split2_merge0_awextras[(EXTRAS - 1):0])
    ,.a_awid(split2_merge0_awid[(IDWID - 1):0])
    ,.a_awlen(split2_merge0_awlen[7:0])
    ,.a_awready(split2_merge0_awready)
    ,.a_awvalid(split2_merge0_awvalid)
    ,.a_bid(split2_merge0_bid[(IDWID - 1):0])
    ,.a_bready(split2_merge0_bready)
    ,.a_bresp(split2_merge0_bresp[1:0])
    ,.a_bvalid(split2_merge0_bvalid)
    ,.a_rdata(split2_merge0_rdata[(DWID - 1):0])
    ,.a_rid(split2_merge0_rid[(IDWID - 1):0])
    ,.a_rlast(split2_merge0_rlast)
    ,.a_rready(split2_merge0_rready)
    ,.a_rresp(split2_merge0_rresp[1:0])
    ,.a_rvalid(split2_merge0_rvalid)
    ,.a_wdata(split2_merge0_wdata[(DWID - 1):0])
    ,.a_wlast(split2_merge0_wlast)
    ,.a_wready(split2_merge0_wready)
    ,.a_wstrb(split2_merge0_wstrb[(WSTRB - 1):0])
    ,.a_wvalid(split2_merge0_wvalid)
    ,.b_araddr(split2_merge1_araddr[31:0])
    ,.b_arburst(split2_merge1_arburst[1:0])
    ,.b_arextras(split2_merge1_arextras[(EXTRAS - 1):0])
    ,.b_arid(split2_merge1_arid[(IDWID - 1):0])
    ,.b_arlen(split2_merge1_arlen[7:0])
    ,.b_arready(split2_merge1_arready)
    ,.b_arvalid(split2_merge1_arvalid)
    ,.b_awaddr(split2_merge1_awaddr[31:0])
    ,.b_awburst(split2_merge1_awburst[1:0])
    ,.b_awextras(split2_merge1_awextras[(EXTRAS - 1):0])
    ,.b_awid(split2_merge1_awid[(IDWID - 1):0])
    ,.b_awlen(split2_merge1_awlen[7:0])
    ,.b_awready(split2_merge1_awready)
    ,.b_awvalid(split2_merge1_awvalid)
    ,.b_bid(split2_merge1_bid[(IDWID - 1):0])
    ,.b_bready(split2_merge1_bready)
    ,.b_bresp(split2_merge1_bresp[1:0])
    ,.b_bvalid(split2_merge1_bvalid)
    ,.b_rdata(split2_merge1_rdata[(DWID - 1):0])
    ,.b_rid(split2_merge1_rid[(IDWID - 1):0])
    ,.b_rlast(split2_merge1_rlast)
    ,.b_rready(split2_merge1_rready)
    ,.b_rresp(split2_merge1_rresp[1:0])
    ,.b_rvalid(split2_merge1_rvalid)
    ,.b_wdata(split2_merge1_wdata[(DWID - 1):0])
    ,.b_wlast(split2_merge1_wlast)
    ,.b_wready(split2_merge1_wready)
    ,.b_wstrb(split2_merge1_wstrb[(WSTRB - 1):0])
    ,.b_wvalid(split2_merge1_wvalid)
    ,.c_araddr(split2_merge2_araddr[31:0])
    ,.c_arburst(split2_merge2_arburst[1:0])
    ,.c_arextras(split2_merge2_arextras[(EXTRAS - 1):0])
    ,.c_arid(split2_merge2_arid[(IDWID - 1):0])
    ,.c_arlen(split2_merge2_arlen[7:0])
    ,.c_arready(split2_merge2_arready)
    ,.c_arvalid(split2_merge2_arvalid)
    ,.c_awaddr(split2_merge2_awaddr[31:0])
    ,.c_awburst(split2_merge2_awburst[1:0])
    ,.c_awextras(split2_merge2_awextras[(EXTRAS - 1):0])
    ,.c_awid(split2_merge2_awid[(IDWID - 1):0])
    ,.c_awlen(split2_merge2_awlen[7:0])
    ,.c_awready(split2_merge2_awready)
    ,.c_awvalid(split2_merge2_awvalid)
    ,.c_bid(split2_merge2_bid[(IDWID - 1):0])
    ,.c_bready(split2_merge2_bready)
    ,.c_bresp(split2_merge2_bresp[1:0])
    ,.c_bvalid(split2_merge2_bvalid)
    ,.c_rdata(split2_merge2_rdata[(DWID - 1):0])
    ,.c_rid(split2_merge2_rid[(IDWID - 1):0])
    ,.c_rlast(split2_merge2_rlast)
    ,.c_rready(split2_merge2_rready)
    ,.c_rresp(split2_merge2_rresp[1:0])
    ,.c_rvalid(split2_merge2_rvalid)
    ,.c_wdata(split2_merge2_wdata[(DWID - 1):0])
    ,.c_wlast(split2_merge2_wlast)
    ,.c_wready(split2_merge2_wready)
    ,.c_wstrb(split2_merge2_wstrb[(WSTRB - 1):0])
    ,.c_wvalid(split2_merge2_wvalid)
    ,.d_araddr(split2_merge3_araddr[31:0])
    ,.d_arburst(split2_merge3_arburst[1:0])
    ,.d_arextras(split2_merge3_arextras[(EXTRAS - 1):0])
    ,.d_arid(split2_merge3_arid[(IDWID - 1):0])
    ,.d_arlen(split2_merge3_arlen[7:0])
    ,.d_arready(split2_merge3_arready)
    ,.d_arvalid(split2_merge3_arvalid)
    ,.d_awaddr(split2_merge3_awaddr[31:0])
    ,.d_awburst(split2_merge3_awburst[1:0])
    ,.d_awextras(split2_merge3_awextras[(EXTRAS - 1):0])
    ,.d_awid(split2_merge3_awid[(IDWID - 1):0])
    ,.d_awlen(split2_merge3_awlen[7:0])
    ,.d_awready(split2_merge3_awready)
    ,.d_awvalid(split2_merge3_awvalid)
    ,.d_bid(split2_merge3_bid[(IDWID - 1):0])
    ,.d_bready(split2_merge3_bready)
    ,.d_bresp(split2_merge3_bresp[1:0])
    ,.d_bvalid(split2_merge3_bvalid)
    ,.d_rdata(split2_merge3_rdata[(DWID - 1):0])
    ,.d_rid(split2_merge3_rid[(IDWID - 1):0])
    ,.d_rlast(split2_merge3_rlast)
    ,.d_rready(split2_merge3_rready)
    ,.d_rresp(split2_merge3_rresp[1:0])
    ,.d_rvalid(split2_merge3_rvalid)
    ,.d_wdata(split2_merge3_wdata[(DWID - 1):0])
    ,.d_wlast(split2_merge3_wlast)
    ,.d_wready(split2_merge3_wready)
    ,.d_wstrb(split2_merge3_wstrb[(WSTRB - 1):0])
    ,.d_wvalid(split2_merge3_wvalid)

);

axi_4_splitter split3 (
     .clk(clk) ,.rst_n(rst_n)

    ,.araddr(mst3_araddr[31:0])
    ,.arburst(mst3_arburst[1:0])
    ,.arextras(mst3_arextras[(EXTRAS - 1):0])
    ,.arid(mst3_arid[(IDWID - 1):0])
    ,.arlen(mst3_arlen[7:0])
    ,.arready(mst3_arready)
    ,.arvalid(mst3_arvalid)
    ,.awaddr(mst3_awaddr[31:0])
    ,.awburst(mst3_awburst[1:0])
    ,.awextras(mst3_awextras[(EXTRAS - 1):0])
    ,.awid(mst3_awid[3:0])
    ,.awlen(mst3_awlen[7:0])
    ,.awready(mst3_awready)
    ,.awvalid(mst3_awvalid)
    ,.bid(mst3_bid[(IDWID - 1):0])
    ,.bready(mst3_bready)
    ,.bresp(mst3_bresp[1:0])
    ,.bvalid(mst3_bvalid)
    ,.rdata(mst3_rdata[(DWID - 1):0])
    ,.rid(mst3_rid[(IDWID - 1):0])
    ,.rlast(mst3_rlast)
    ,.rready(mst3_rready)
    ,.rresp(mst3_rresp[1:0])
    ,.rvalid(mst3_rvalid)
    ,.wdata(mst3_wdata[(DWID - 1):0])
    ,.wlast(mst3_wlast)
    ,.wready(mst3_wready)
    ,.wstrb(mst3_wstrb[(WSTRB - 1):0])
    ,.wvalid(mst3_wvalid)

    ,.a_araddr(split3_merge0_araddr[31:0])
    ,.a_arburst(split3_merge0_arburst[1:0])
    ,.a_arextras(split3_merge0_arextras[(EXTRAS - 1):0])
    ,.a_arid(split3_merge0_arid[(IDWID - 1):0])
    ,.a_arlen(split3_merge0_arlen[7:0])
    ,.a_arready(split3_merge0_arready)
    ,.a_arvalid(split3_merge0_arvalid)
    ,.a_awaddr(split3_merge0_awaddr[31:0])
    ,.a_awburst(split3_merge0_awburst[1:0])
    ,.a_awextras(split3_merge0_awextras[(EXTRAS - 1):0])
    ,.a_awid(split3_merge0_awid[(IDWID - 1):0])
    ,.a_awlen(split3_merge0_awlen[7:0])
    ,.a_awready(split3_merge0_awready)
    ,.a_awvalid(split3_merge0_awvalid)
    ,.a_bid(split3_merge0_bid[(IDWID - 1):0])
    ,.a_bready(split3_merge0_bready)
    ,.a_bresp(split3_merge0_bresp[1:0])
    ,.a_bvalid(split3_merge0_bvalid)
    ,.a_rdata(split3_merge0_rdata[(DWID - 1):0])
    ,.a_rid(split3_merge0_rid[(IDWID - 1):0])
    ,.a_rlast(split3_merge0_rlast)
    ,.a_rready(split3_merge0_rready)
    ,.a_rresp(split3_merge0_rresp[1:0])
    ,.a_rvalid(split3_merge0_rvalid)
    ,.a_wdata(split3_merge0_wdata[(DWID - 1):0])
    ,.a_wlast(split3_merge0_wlast)
    ,.a_wready(split3_merge0_wready)
    ,.a_wstrb(split3_merge0_wstrb[(WSTRB - 1):0])
    ,.a_wvalid(split3_merge0_wvalid)
    ,.b_araddr(split3_merge1_araddr[31:0])
    ,.b_arburst(split3_merge1_arburst[1:0])
    ,.b_arextras(split3_merge1_arextras[(EXTRAS - 1):0])
    ,.b_arid(split3_merge1_arid[(IDWID - 1):0])
    ,.b_arlen(split3_merge1_arlen[7:0])
    ,.b_arready(split3_merge1_arready)
    ,.b_arvalid(split3_merge1_arvalid)
    ,.b_awaddr(split3_merge1_awaddr[31:0])
    ,.b_awburst(split3_merge1_awburst[1:0])
    ,.b_awextras(split3_merge1_awextras[(EXTRAS - 1):0])
    ,.b_awid(split3_merge1_awid[(IDWID - 1):0])
    ,.b_awlen(split3_merge1_awlen[7:0])
    ,.b_awready(split3_merge1_awready)
    ,.b_awvalid(split3_merge1_awvalid)
    ,.b_bid(split3_merge1_bid[(IDWID - 1):0])
    ,.b_bready(split3_merge1_bready)
    ,.b_bresp(split3_merge1_bresp[1:0])
    ,.b_bvalid(split3_merge1_bvalid)
    ,.b_rdata(split3_merge1_rdata[(DWID - 1):0])
    ,.b_rid(split3_merge1_rid[(IDWID - 1):0])
    ,.b_rlast(split3_merge1_rlast)
    ,.b_rready(split3_merge1_rready)
    ,.b_rresp(split3_merge1_rresp[1:0])
    ,.b_rvalid(split3_merge1_rvalid)
    ,.b_wdata(split3_merge1_wdata[(DWID - 1):0])
    ,.b_wlast(split3_merge1_wlast)
    ,.b_wready(split3_merge1_wready)
    ,.b_wstrb(split3_merge1_wstrb[(WSTRB - 1):0])
    ,.b_wvalid(split3_merge1_wvalid)
    ,.c_araddr(split3_merge2_araddr[31:0])
    ,.c_arburst(split3_merge2_arburst[1:0])
    ,.c_arextras(split3_merge2_arextras[(EXTRAS - 1):0])
    ,.c_arid(split3_merge2_arid[(IDWID - 1):0])
    ,.c_arlen(split3_merge2_arlen[7:0])
    ,.c_arready(split3_merge2_arready)
    ,.c_arvalid(split3_merge2_arvalid)
    ,.c_awaddr(split3_merge2_awaddr[31:0])
    ,.c_awburst(split3_merge2_awburst[1:0])
    ,.c_awextras(split3_merge2_awextras[(EXTRAS - 1):0])
    ,.c_awid(split3_merge2_awid[(IDWID - 1):0])
    ,.c_awlen(split3_merge2_awlen[7:0])
    ,.c_awready(split3_merge2_awready)
    ,.c_awvalid(split3_merge2_awvalid)
    ,.c_bid(split3_merge2_bid[(IDWID - 1):0])
    ,.c_bready(split3_merge2_bready)
    ,.c_bresp(split3_merge2_bresp[1:0])
    ,.c_bvalid(split3_merge2_bvalid)
    ,.c_rdata(split3_merge2_rdata[(DWID - 1):0])
    ,.c_rid(split3_merge2_rid[(IDWID - 1):0])
    ,.c_rlast(split3_merge2_rlast)
    ,.c_rready(split3_merge2_rready)
    ,.c_rresp(split3_merge2_rresp[1:0])
    ,.c_rvalid(split3_merge2_rvalid)
    ,.c_wdata(split3_merge2_wdata[(DWID - 1):0])
    ,.c_wlast(split3_merge2_wlast)
    ,.c_wready(split3_merge2_wready)
    ,.c_wstrb(split3_merge2_wstrb[(WSTRB - 1):0])
    ,.c_wvalid(split3_merge2_wvalid)
    ,.d_araddr(split3_merge3_araddr[31:0])
    ,.d_arburst(split3_merge3_arburst[1:0])
    ,.d_arextras(split3_merge3_arextras[(EXTRAS - 1):0])
    ,.d_arid(split3_merge3_arid[(IDWID - 1):0])
    ,.d_arlen(split3_merge3_arlen[7:0])
    ,.d_arready(split3_merge3_arready)
    ,.d_arvalid(split3_merge3_arvalid)
    ,.d_awaddr(split3_merge3_awaddr[31:0])
    ,.d_awburst(split3_merge3_awburst[1:0])
    ,.d_awextras(split3_merge3_awextras[(EXTRAS - 1):0])
    ,.d_awid(split3_merge3_awid[(IDWID - 1):0])
    ,.d_awlen(split3_merge3_awlen[7:0])
    ,.d_awready(split3_merge3_awready)
    ,.d_awvalid(split3_merge3_awvalid)
    ,.d_bid(split3_merge3_bid[(IDWID - 1):0])
    ,.d_bready(split3_merge3_bready)
    ,.d_bresp(split3_merge3_bresp[1:0])
    ,.d_bvalid(split3_merge3_bvalid)
    ,.d_rdata(split3_merge3_rdata[(DWID - 1):0])
    ,.d_rid(split3_merge3_rid[(IDWID - 1):0])
    ,.d_rlast(split3_merge3_rlast)
    ,.d_rready(split3_merge3_rready)
    ,.d_rresp(split3_merge3_rresp[1:0])
    ,.d_rvalid(split3_merge3_rvalid)
    ,.d_wdata(split3_merge3_wdata[(DWID - 1):0])
    ,.d_wlast(split3_merge3_wlast)
    ,.d_wready(split3_merge3_wready)
    ,.d_wstrb(split3_merge3_wstrb[(WSTRB - 1):0])
    ,.d_wvalid(split3_merge3_wvalid)

);

wire [IDWID-1:0] split4_merge4_arid ;
wire [31:0] split4_merge4_araddr ;
wire [7:0] split4_merge4_arlen ;
wire [EXTRAS-1:0] split4_merge4_arextras ;
wire [1:0] split4_merge4_arburst ;
wire split4_merge4_arvalid ;
wire split4_merge4_arready ;
wire [IDWID-1:0] split4_merge4_rid ;
wire [DWID-1:0] split4_merge4_rdata ;
wire [1:0] split4_merge4_rresp ;
wire split4_merge4_rlast ;
wire split4_merge4_rvalid ;
wire split4_merge4_rready ;

wire [IDWID-1:0] split4_merge4_awid ;
wire [31:0] split4_merge4_awaddr ;
wire [7:0] split4_merge4_awlen ;
wire [EXTRAS-1:0] split4_merge4_awextras ;
wire [1:0] split4_merge4_awburst ;
wire split4_merge4_awvalid ;
wire split4_merge4_awready ;
wire [DWID-1:0] split4_merge4_wdata ;
wire [WSTRB-1:0] split4_merge4_wstrb ;
wire split4_merge4_wlast ;
wire split4_merge4_wvalid ;
wire split4_merge4_wready ;
wire [IDWID-1:0] split4_merge4_bid ;
wire [1:0] split4_merge4_bresp ;
wire split4_merge4_bvalid ;
wire split4_merge4_bready ;


wire [IDWID-1:0] split4_merge5_arid ;
wire [31:0] split4_merge5_araddr ;
wire [7:0] split4_merge5_arlen ;
wire [EXTRAS-1:0] split4_merge5_arextras ;
wire [1:0] split4_merge5_arburst ;
wire split4_merge5_arvalid ;
wire split4_merge5_arready ;
wire [IDWID-1:0] split4_merge5_rid ;
wire [DWID-1:0] split4_merge5_rdata ;
wire [1:0] split4_merge5_rresp ;
wire split4_merge5_rlast ;
wire split4_merge5_rvalid ;
wire split4_merge5_rready ;

wire [IDWID-1:0] split4_merge5_awid ;
wire [31:0] split4_merge5_awaddr ;
wire [7:0] split4_merge5_awlen ;
wire [EXTRAS-1:0] split4_merge5_awextras ;
wire [1:0] split4_merge5_awburst ;
wire split4_merge5_awvalid ;
wire split4_merge5_awready ;
wire [DWID-1:0] split4_merge5_wdata ;
wire [WSTRB-1:0] split4_merge5_wstrb ;
wire split4_merge5_wlast ;
wire split4_merge5_wvalid ;
wire split4_merge5_wready ;
wire [IDWID-1:0] split4_merge5_bid ;
wire [1:0] split4_merge5_bresp ;
wire split4_merge5_bvalid ;
wire split4_merge5_bready ;


wire [IDWID-1:0] split4_merge6_arid ;
wire [31:0] split4_merge6_araddr ;
wire [7:0] split4_merge6_arlen ;
wire [EXTRAS-1:0] split4_merge6_arextras ;
wire [1:0] split4_merge6_arburst ;
wire split4_merge6_arvalid ;
wire split4_merge6_arready ;
wire [IDWID-1:0] split4_merge6_rid ;
wire [DWID-1:0] split4_merge6_rdata ;
wire [1:0] split4_merge6_rresp ;
wire split4_merge6_rlast ;
wire split4_merge6_rvalid ;
wire split4_merge6_rready ;

wire [IDWID-1:0] split4_merge6_awid ;
wire [31:0] split4_merge6_awaddr ;
wire [7:0] split4_merge6_awlen ;
wire [EXTRAS-1:0] split4_merge6_awextras ;
wire [1:0] split4_merge6_awburst ;
wire split4_merge6_awvalid ;
wire split4_merge6_awready ;
wire [DWID-1:0] split4_merge6_wdata ;
wire [WSTRB-1:0] split4_merge6_wstrb ;
wire split4_merge6_wlast ;
wire split4_merge6_wvalid ;
wire split4_merge6_wready ;
wire [IDWID-1:0] split4_merge6_bid ;
wire [1:0] split4_merge6_bresp ;
wire split4_merge6_bvalid ;
wire split4_merge6_bready ;


wire [IDWID-1:0] split4_merge7_arid ;
wire [31:0] split4_merge7_araddr ;
wire [7:0] split4_merge7_arlen ;
wire [EXTRAS-1:0] split4_merge7_arextras ;
wire [1:0] split4_merge7_arburst ;
wire split4_merge7_arvalid ;
wire split4_merge7_arready ;
wire [IDWID-1:0] split4_merge7_rid ;
wire [DWID-1:0] split4_merge7_rdata ;
wire [1:0] split4_merge7_rresp ;
wire split4_merge7_rlast ;
wire split4_merge7_rvalid ;
wire split4_merge7_rready ;

wire [IDWID-1:0] split4_merge7_awid ;
wire [31:0] split4_merge7_awaddr ;
wire [7:0] split4_merge7_awlen ;
wire [EXTRAS-1:0] split4_merge7_awextras ;
wire [1:0] split4_merge7_awburst ;
wire split4_merge7_awvalid ;
wire split4_merge7_awready ;
wire [DWID-1:0] split4_merge7_wdata ;
wire [WSTRB-1:0] split4_merge7_wstrb ;
wire split4_merge7_wlast ;
wire split4_merge7_wvalid ;
wire split4_merge7_wready ;
wire [IDWID-1:0] split4_merge7_bid ;
wire [1:0] split4_merge7_bresp ;
wire split4_merge7_bvalid ;
wire split4_merge7_bready ;


axi_4_splitter split4 (
     .clk(clk) ,.rst_n(rst_n)

    ,.araddr(mst4_araddr[31:0])
    ,.arburst(mst4_arburst[1:0])
    ,.arextras(mst4_arextras[(EXTRAS - 1):0])
    ,.arid(mst4_arid[(IDWID - 1):0])
    ,.arlen(mst4_arlen[7:0])
    ,.arready(mst4_arready)
    ,.arvalid(mst4_arvalid)
    ,.awaddr(mst4_awaddr[31:0])
    ,.awburst(mst4_awburst[1:0])
    ,.awextras(mst4_awextras[(EXTRAS - 1):0])
    ,.awid(mst4_awid[3:0])
    ,.awlen(mst4_awlen[7:0])
    ,.awready(mst4_awready)
    ,.awvalid(mst4_awvalid)
    ,.bid(mst4_bid[(IDWID - 1):0])
    ,.bready(mst4_bready)
    ,.bresp(mst4_bresp[1:0])
    ,.bvalid(mst4_bvalid)
    ,.rdata(mst4_rdata[(DWID - 1):0])
    ,.rid(mst4_rid[(IDWID - 1):0])
    ,.rlast(mst4_rlast)
    ,.rready(mst4_rready)
    ,.rresp(mst4_rresp[1:0])
    ,.rvalid(mst4_rvalid)
    ,.wdata(mst4_wdata[(DWID - 1):0])
    ,.wlast(mst4_wlast)
    ,.wready(mst4_wready)
    ,.wstrb(mst4_wstrb[(WSTRB - 1):0])
    ,.wvalid(mst4_wvalid)

    ,.a_araddr(split4_merge4_araddr[31:0])
    ,.a_arburst(split4_merge4_arburst[1:0])
    ,.a_arextras(split4_merge4_arextras[(EXTRAS - 1):0])
    ,.a_arid(split4_merge4_arid[(IDWID - 1):0])
    ,.a_arlen(split4_merge4_arlen[7:0])
    ,.a_arready(split4_merge4_arready)
    ,.a_arvalid(split4_merge4_arvalid)
    ,.a_awaddr(split4_merge4_awaddr[31:0])
    ,.a_awburst(split4_merge4_awburst[1:0])
    ,.a_awextras(split4_merge4_awextras[(EXTRAS - 1):0])
    ,.a_awid(split4_merge4_awid[(IDWID - 1):0])
    ,.a_awlen(split4_merge4_awlen[7:0])
    ,.a_awready(split4_merge4_awready)
    ,.a_awvalid(split4_merge4_awvalid)
    ,.a_bid(split4_merge4_bid[(IDWID - 1):0])
    ,.a_bready(split4_merge4_bready)
    ,.a_bresp(split4_merge4_bresp[1:0])
    ,.a_bvalid(split4_merge4_bvalid)
    ,.a_rdata(split4_merge4_rdata[(DWID - 1):0])
    ,.a_rid(split4_merge4_rid[(IDWID - 1):0])
    ,.a_rlast(split4_merge4_rlast)
    ,.a_rready(split4_merge4_rready)
    ,.a_rresp(split4_merge4_rresp[1:0])
    ,.a_rvalid(split4_merge4_rvalid)
    ,.a_wdata(split4_merge4_wdata[(DWID - 1):0])
    ,.a_wlast(split4_merge4_wlast)
    ,.a_wready(split4_merge4_wready)
    ,.a_wstrb(split4_merge4_wstrb[(WSTRB - 1):0])
    ,.a_wvalid(split4_merge4_wvalid)
    ,.b_araddr(split4_merge5_araddr[31:0])
    ,.b_arburst(split4_merge5_arburst[1:0])
    ,.b_arextras(split4_merge5_arextras[(EXTRAS - 1):0])
    ,.b_arid(split4_merge5_arid[(IDWID - 1):0])
    ,.b_arlen(split4_merge5_arlen[7:0])
    ,.b_arready(split4_merge5_arready)
    ,.b_arvalid(split4_merge5_arvalid)
    ,.b_awaddr(split4_merge5_awaddr[31:0])
    ,.b_awburst(split4_merge5_awburst[1:0])
    ,.b_awextras(split4_merge5_awextras[(EXTRAS - 1):0])
    ,.b_awid(split4_merge5_awid[(IDWID - 1):0])
    ,.b_awlen(split4_merge5_awlen[7:0])
    ,.b_awready(split4_merge5_awready)
    ,.b_awvalid(split4_merge5_awvalid)
    ,.b_bid(split4_merge5_bid[(IDWID - 1):0])
    ,.b_bready(split4_merge5_bready)
    ,.b_bresp(split4_merge5_bresp[1:0])
    ,.b_bvalid(split4_merge5_bvalid)
    ,.b_rdata(split4_merge5_rdata[(DWID - 1):0])
    ,.b_rid(split4_merge5_rid[(IDWID - 1):0])
    ,.b_rlast(split4_merge5_rlast)
    ,.b_rready(split4_merge5_rready)
    ,.b_rresp(split4_merge5_rresp[1:0])
    ,.b_rvalid(split4_merge5_rvalid)
    ,.b_wdata(split4_merge5_wdata[(DWID - 1):0])
    ,.b_wlast(split4_merge5_wlast)
    ,.b_wready(split4_merge5_wready)
    ,.b_wstrb(split4_merge5_wstrb[(WSTRB - 1):0])
    ,.b_wvalid(split4_merge5_wvalid)
    ,.c_araddr(split4_merge6_araddr[31:0])
    ,.c_arburst(split4_merge6_arburst[1:0])
    ,.c_arextras(split4_merge6_arextras[(EXTRAS - 1):0])
    ,.c_arid(split4_merge6_arid[(IDWID - 1):0])
    ,.c_arlen(split4_merge6_arlen[7:0])
    ,.c_arready(split4_merge6_arready)
    ,.c_arvalid(split4_merge6_arvalid)
    ,.c_awaddr(split4_merge6_awaddr[31:0])
    ,.c_awburst(split4_merge6_awburst[1:0])
    ,.c_awextras(split4_merge6_awextras[(EXTRAS - 1):0])
    ,.c_awid(split4_merge6_awid[(IDWID - 1):0])
    ,.c_awlen(split4_merge6_awlen[7:0])
    ,.c_awready(split4_merge6_awready)
    ,.c_awvalid(split4_merge6_awvalid)
    ,.c_bid(split4_merge6_bid[(IDWID - 1):0])
    ,.c_bready(split4_merge6_bready)
    ,.c_bresp(split4_merge6_bresp[1:0])
    ,.c_bvalid(split4_merge6_bvalid)
    ,.c_rdata(split4_merge6_rdata[(DWID - 1):0])
    ,.c_rid(split4_merge6_rid[(IDWID - 1):0])
    ,.c_rlast(split4_merge6_rlast)
    ,.c_rready(split4_merge6_rready)
    ,.c_rresp(split4_merge6_rresp[1:0])
    ,.c_rvalid(split4_merge6_rvalid)
    ,.c_wdata(split4_merge6_wdata[(DWID - 1):0])
    ,.c_wlast(split4_merge6_wlast)
    ,.c_wready(split4_merge6_wready)
    ,.c_wstrb(split4_merge6_wstrb[(WSTRB - 1):0])
    ,.c_wvalid(split4_merge6_wvalid)
    ,.d_araddr(split4_merge7_araddr[31:0])
    ,.d_arburst(split4_merge7_arburst[1:0])
    ,.d_arextras(split4_merge7_arextras[(EXTRAS - 1):0])
    ,.d_arid(split4_merge7_arid[(IDWID - 1):0])
    ,.d_arlen(split4_merge7_arlen[7:0])
    ,.d_arready(split4_merge7_arready)
    ,.d_arvalid(split4_merge7_arvalid)
    ,.d_awaddr(split4_merge7_awaddr[31:0])
    ,.d_awburst(split4_merge7_awburst[1:0])
    ,.d_awextras(split4_merge7_awextras[(EXTRAS - 1):0])
    ,.d_awid(split4_merge7_awid[(IDWID - 1):0])
    ,.d_awlen(split4_merge7_awlen[7:0])
    ,.d_awready(split4_merge7_awready)
    ,.d_awvalid(split4_merge7_awvalid)
    ,.d_bid(split4_merge7_bid[(IDWID - 1):0])
    ,.d_bready(split4_merge7_bready)
    ,.d_bresp(split4_merge7_bresp[1:0])
    ,.d_bvalid(split4_merge7_bvalid)
    ,.d_rdata(split4_merge7_rdata[(DWID - 1):0])
    ,.d_rid(split4_merge7_rid[(IDWID - 1):0])
    ,.d_rlast(split4_merge7_rlast)
    ,.d_rready(split4_merge7_rready)
    ,.d_rresp(split4_merge7_rresp[1:0])
    ,.d_rvalid(split4_merge7_rvalid)
    ,.d_wdata(split4_merge7_wdata[(DWID - 1):0])
    ,.d_wlast(split4_merge7_wlast)
    ,.d_wready(split4_merge7_wready)
    ,.d_wstrb(split4_merge7_wstrb[(WSTRB - 1):0])
    ,.d_wvalid(split4_merge7_wvalid)

);

wire [IDWID-1:0] merge4_split104_arid ;
wire [31:0] merge4_split104_araddr ;
wire [7:0] merge4_split104_arlen ;
wire [EXTRAS-1:0] merge4_split104_arextras ;
wire [1:0] merge4_split104_arburst ;
wire merge4_split104_arvalid ;
wire merge4_split104_arready ;
wire [IDWID-1:0] merge4_split104_rid ;
wire [DWID-1:0] merge4_split104_rdata ;
wire [1:0] merge4_split104_rresp ;
wire merge4_split104_rlast ;
wire merge4_split104_rvalid ;
wire merge4_split104_rready ;

wire [IDWID-1:0] merge4_split104_awid ;
wire [31:0] merge4_split104_awaddr ;
wire [7:0] merge4_split104_awlen ;
wire [EXTRAS-1:0] merge4_split104_awextras ;
wire [1:0] merge4_split104_awburst ;
wire merge4_split104_awvalid ;
wire merge4_split104_awready ;
wire [DWID-1:0] merge4_split104_wdata ;
wire [WSTRB-1:0] merge4_split104_wstrb ;
wire merge4_split104_wlast ;
wire merge4_split104_wvalid ;
wire merge4_split104_wready ;
wire [IDWID-1:0] merge4_split104_bid ;
wire [1:0] merge4_split104_bresp ;
wire merge4_split104_bvalid ;
wire merge4_split104_bready ;


wire [IDWID-1:0] split5_merge4_arid ;
wire [31:0] split5_merge4_araddr ;
wire [7:0] split5_merge4_arlen ;
wire [EXTRAS-1:0] split5_merge4_arextras ;
wire [1:0] split5_merge4_arburst ;
wire split5_merge4_arvalid ;
wire split5_merge4_arready ;
wire [IDWID-1:0] split5_merge4_rid ;
wire [DWID-1:0] split5_merge4_rdata ;
wire [1:0] split5_merge4_rresp ;
wire split5_merge4_rlast ;
wire split5_merge4_rvalid ;
wire split5_merge4_rready ;

wire [IDWID-1:0] split5_merge4_awid ;
wire [31:0] split5_merge4_awaddr ;
wire [7:0] split5_merge4_awlen ;
wire [EXTRAS-1:0] split5_merge4_awextras ;
wire [1:0] split5_merge4_awburst ;
wire split5_merge4_awvalid ;
wire split5_merge4_awready ;
wire [DWID-1:0] split5_merge4_wdata ;
wire [WSTRB-1:0] split5_merge4_wstrb ;
wire split5_merge4_wlast ;
wire split5_merge4_wvalid ;
wire split5_merge4_wready ;
wire [IDWID-1:0] split5_merge4_bid ;
wire [1:0] split5_merge4_bresp ;
wire split5_merge4_bvalid ;
wire split5_merge4_bready ;


wire [IDWID-1:0] split6_merge4_arid ;
wire [31:0] split6_merge4_araddr ;
wire [7:0] split6_merge4_arlen ;
wire [EXTRAS-1:0] split6_merge4_arextras ;
wire [1:0] split6_merge4_arburst ;
wire split6_merge4_arvalid ;
wire split6_merge4_arready ;
wire [IDWID-1:0] split6_merge4_rid ;
wire [DWID-1:0] split6_merge4_rdata ;
wire [1:0] split6_merge4_rresp ;
wire split6_merge4_rlast ;
wire split6_merge4_rvalid ;
wire split6_merge4_rready ;

wire [IDWID-1:0] split6_merge4_awid ;
wire [31:0] split6_merge4_awaddr ;
wire [7:0] split6_merge4_awlen ;
wire [EXTRAS-1:0] split6_merge4_awextras ;
wire [1:0] split6_merge4_awburst ;
wire split6_merge4_awvalid ;
wire split6_merge4_awready ;
wire [DWID-1:0] split6_merge4_wdata ;
wire [WSTRB-1:0] split6_merge4_wstrb ;
wire split6_merge4_wlast ;
wire split6_merge4_wvalid ;
wire split6_merge4_wready ;
wire [IDWID-1:0] split6_merge4_bid ;
wire [1:0] split6_merge4_bresp ;
wire split6_merge4_bvalid ;
wire split6_merge4_bready ;


wire [IDWID-1:0] split7_merge4_arid ;
wire [31:0] split7_merge4_araddr ;
wire [7:0] split7_merge4_arlen ;
wire [EXTRAS-1:0] split7_merge4_arextras ;
wire [1:0] split7_merge4_arburst ;
wire split7_merge4_arvalid ;
wire split7_merge4_arready ;
wire [IDWID-1:0] split7_merge4_rid ;
wire [DWID-1:0] split7_merge4_rdata ;
wire [1:0] split7_merge4_rresp ;
wire split7_merge4_rlast ;
wire split7_merge4_rvalid ;
wire split7_merge4_rready ;

wire [IDWID-1:0] split7_merge4_awid ;
wire [31:0] split7_merge4_awaddr ;
wire [7:0] split7_merge4_awlen ;
wire [EXTRAS-1:0] split7_merge4_awextras ;
wire [1:0] split7_merge4_awburst ;
wire split7_merge4_awvalid ;
wire split7_merge4_awready ;
wire [DWID-1:0] split7_merge4_wdata ;
wire [WSTRB-1:0] split7_merge4_wstrb ;
wire split7_merge4_wlast ;
wire split7_merge4_wvalid ;
wire split7_merge4_wready ;
wire [IDWID-1:0] split7_merge4_bid ;
wire [1:0] split7_merge4_bresp ;
wire split7_merge4_bvalid ;
wire split7_merge4_bready ;


axi_4_merger merge4 (
     .clk(clk),.rst_n(rst_n)
    ,.araddr(merge4_split104_araddr[31:0])
    ,.arburst(merge4_split104_arburst[1:0])
    ,.arextras(merge4_split104_arextras[(EXTRAS - 1):0])
    ,.arid(merge4_split104_arid[(IDWID - 1):0])
    ,.arlen(merge4_split104_arlen[7:0])
    ,.arready(merge4_split104_arready)
    ,.arvalid(merge4_split104_arvalid)
    ,.awaddr(merge4_split104_awaddr[31:0])
    ,.awburst(merge4_split104_awburst[1:0])
    ,.awextras(merge4_split104_awextras[(EXTRAS - 1):0])
    ,.awid(merge4_split104_awid[3:0])
    ,.awlen(merge4_split104_awlen[7:0])
    ,.awready(merge4_split104_awready)
    ,.awvalid(merge4_split104_awvalid)
    ,.bid(merge4_split104_bid[(IDWID - 1):0])
    ,.bready(merge4_split104_bready)
    ,.bresp(merge4_split104_bresp[1:0])
    ,.bvalid(merge4_split104_bvalid)
    ,.rid(merge4_split104_rid[(IDWID - 1):0])
    ,.rlast(merge4_split104_rlast)
    ,.rready(merge4_split104_rready)
    ,.rresp(merge4_split104_rresp[1:0])
    ,.rvalid(merge4_split104_rvalid)
    ,.rdata(merge4_split104_rdata[(DWID - 1):0])
    ,.wdata(merge4_split104_wdata[(DWID - 1):0])
    ,.wlast(merge4_split104_wlast)
    ,.wready(merge4_split104_wready)
    ,.wstrb(merge4_split104_wstrb[(WSTRB - 1):0])
    ,.wvalid(merge4_split104_wvalid)


    ,.a_araddr(split4_merge4_araddr[31:0])
    ,.a_arburst(split4_merge4_arburst[1:0])
    ,.a_arextras(split4_merge4_arextras[(EXTRAS - 1):0])
    ,.a_arid(split4_merge4_arid[(IDWID - 1):0])
    ,.a_arlen(split4_merge4_arlen[7:0])
    ,.a_arready(split4_merge4_arready)
    ,.a_arvalid(split4_merge4_arvalid)
    ,.a_awaddr(split4_merge4_awaddr[31:0])
    ,.a_awburst(split4_merge4_awburst[1:0])
    ,.a_awextras(split4_merge4_awextras[(EXTRAS - 1):0])
    ,.a_awid(split4_merge4_awid[(IDWID - 1):0])
    ,.a_awlen(split4_merge4_awlen[7:0])
    ,.a_awready(split4_merge4_awready)
    ,.a_awvalid(split4_merge4_awvalid)
    ,.a_bid(split4_merge4_bid[(IDWID - 1):0])
    ,.a_bready(split4_merge4_bready)
    ,.a_bresp(split4_merge4_bresp[1:0])
    ,.a_bvalid(split4_merge4_bvalid)
    ,.a_rdata(split4_merge4_rdata[(DWID - 1):0])
    ,.a_rid(split4_merge4_rid[(IDWID - 1):0])
    ,.a_rlast(split4_merge4_rlast)
    ,.a_rready(split4_merge4_rready)
    ,.a_rresp(split4_merge4_rresp[1:0])
    ,.a_rvalid(split4_merge4_rvalid)
    ,.a_wdata(split4_merge4_wdata[(DWID - 1):0])
    ,.a_wlast(split4_merge4_wlast)
    ,.a_wready(split4_merge4_wready)
    ,.a_wstrb(split4_merge4_wstrb[(WSTRB - 1):0])
    ,.a_wvalid(split4_merge4_wvalid)

    ,.b_araddr(split5_merge4_araddr[31:0])
    ,.b_arburst(split5_merge4_arburst[1:0])
    ,.b_arextras(split5_merge4_arextras[(EXTRAS - 1):0])
    ,.b_arid(split5_merge4_arid[(IDWID - 1):0])
    ,.b_arlen(split5_merge4_arlen[7:0])
    ,.b_arready(split5_merge4_arready)
    ,.b_arvalid(split5_merge4_arvalid)
    ,.b_awaddr(split5_merge4_awaddr[31:0])
    ,.b_awburst(split5_merge4_awburst[1:0])
    ,.b_awextras(split5_merge4_awextras[(EXTRAS - 1):0])
    ,.b_awid(split5_merge4_awid[(IDWID - 1):0])
    ,.b_awlen(split5_merge4_awlen[7:0])
    ,.b_awready(split5_merge4_awready)
    ,.b_awvalid(split5_merge4_awvalid)
    ,.b_bid(split5_merge4_bid[(IDWID - 1):0])
    ,.b_bready(split5_merge4_bready)
    ,.b_bresp(split5_merge4_bresp[1:0])
    ,.b_bvalid(split5_merge4_bvalid)
    ,.b_rdata(split5_merge4_rdata[(DWID - 1):0])
    ,.b_rid(split5_merge4_rid[(IDWID - 1):0])
    ,.b_rlast(split5_merge4_rlast)
    ,.b_rready(split5_merge4_rready)
    ,.b_rresp(split5_merge4_rresp[1:0])
    ,.b_rvalid(split5_merge4_rvalid)
    ,.b_wdata(split5_merge4_wdata[(DWID - 1):0])
    ,.b_wlast(split5_merge4_wlast)
    ,.b_wready(split5_merge4_wready)
    ,.b_wstrb(split5_merge4_wstrb[(WSTRB - 1):0])
    ,.b_wvalid(split5_merge4_wvalid)

    ,.c_araddr(split6_merge4_araddr[31:0])
    ,.c_arburst(split6_merge4_arburst[1:0])
    ,.c_arextras(split6_merge4_arextras[(EXTRAS - 1):0])
    ,.c_arid(split6_merge4_arid[(IDWID - 1):0])
    ,.c_arlen(split6_merge4_arlen[7:0])
    ,.c_arready(split6_merge4_arready)
    ,.c_arvalid(split6_merge4_arvalid)
    ,.c_awaddr(split6_merge4_awaddr[31:0])
    ,.c_awburst(split6_merge4_awburst[1:0])
    ,.c_awextras(split6_merge4_awextras[(EXTRAS - 1):0])
    ,.c_awid(split6_merge4_awid[(IDWID - 1):0])
    ,.c_awlen(split6_merge4_awlen[7:0])
    ,.c_awready(split6_merge4_awready)
    ,.c_awvalid(split6_merge4_awvalid)
    ,.c_bid(split6_merge4_bid[(IDWID - 1):0])
    ,.c_bready(split6_merge4_bready)
    ,.c_bresp(split6_merge4_bresp[1:0])
    ,.c_bvalid(split6_merge4_bvalid)
    ,.c_rdata(split6_merge4_rdata[(DWID - 1):0])
    ,.c_rid(split6_merge4_rid[(IDWID - 1):0])
    ,.c_rlast(split6_merge4_rlast)
    ,.c_rready(split6_merge4_rready)
    ,.c_rresp(split6_merge4_rresp[1:0])
    ,.c_rvalid(split6_merge4_rvalid)
    ,.c_wdata(split6_merge4_wdata[(DWID - 1):0])
    ,.c_wlast(split6_merge4_wlast)
    ,.c_wready(split6_merge4_wready)
    ,.c_wstrb(split6_merge4_wstrb[(WSTRB - 1):0])
    ,.c_wvalid(split6_merge4_wvalid)

    ,.d_araddr(split7_merge4_araddr[31:0])
    ,.d_arburst(split7_merge4_arburst[1:0])
    ,.d_arextras(split7_merge4_arextras[(EXTRAS - 1):0])
    ,.d_arid(split7_merge4_arid[(IDWID - 1):0])
    ,.d_arlen(split7_merge4_arlen[7:0])
    ,.d_arready(split7_merge4_arready)
    ,.d_arvalid(split7_merge4_arvalid)
    ,.d_awaddr(split7_merge4_awaddr[31:0])
    ,.d_awburst(split7_merge4_awburst[1:0])
    ,.d_awextras(split7_merge4_awextras[(EXTRAS - 1):0])
    ,.d_awid(split7_merge4_awid[(IDWID - 1):0])
    ,.d_awlen(split7_merge4_awlen[7:0])
    ,.d_awready(split7_merge4_awready)
    ,.d_awvalid(split7_merge4_awvalid)
    ,.d_bid(split7_merge4_bid[(IDWID - 1):0])
    ,.d_bready(split7_merge4_bready)
    ,.d_bresp(split7_merge4_bresp[1:0])
    ,.d_bvalid(split7_merge4_bvalid)
    ,.d_rdata(split7_merge4_rdata[(DWID - 1):0])
    ,.d_rid(split7_merge4_rid[(IDWID - 1):0])
    ,.d_rlast(split7_merge4_rlast)
    ,.d_rready(split7_merge4_rready)
    ,.d_rresp(split7_merge4_rresp[1:0])
    ,.d_rvalid(split7_merge4_rvalid)
    ,.d_wdata(split7_merge4_wdata[(DWID - 1):0])
    ,.d_wlast(split7_merge4_wlast)
    ,.d_wready(split7_merge4_wready)
    ,.d_wstrb(split7_merge4_wstrb[(WSTRB - 1):0])
    ,.d_wvalid(split7_merge4_wvalid)
);


wire [IDWID-1:0] merge5_split105_arid ;
wire [31:0] merge5_split105_araddr ;
wire [7:0] merge5_split105_arlen ;
wire [EXTRAS-1:0] merge5_split105_arextras ;
wire [1:0] merge5_split105_arburst ;
wire merge5_split105_arvalid ;
wire merge5_split105_arready ;
wire [IDWID-1:0] merge5_split105_rid ;
wire [DWID-1:0] merge5_split105_rdata ;
wire [1:0] merge5_split105_rresp ;
wire merge5_split105_rlast ;
wire merge5_split105_rvalid ;
wire merge5_split105_rready ;

wire [IDWID-1:0] merge5_split105_awid ;
wire [31:0] merge5_split105_awaddr ;
wire [7:0] merge5_split105_awlen ;
wire [EXTRAS-1:0] merge5_split105_awextras ;
wire [1:0] merge5_split105_awburst ;
wire merge5_split105_awvalid ;
wire merge5_split105_awready ;
wire [DWID-1:0] merge5_split105_wdata ;
wire [WSTRB-1:0] merge5_split105_wstrb ;
wire merge5_split105_wlast ;
wire merge5_split105_wvalid ;
wire merge5_split105_wready ;
wire [IDWID-1:0] merge5_split105_bid ;
wire [1:0] merge5_split105_bresp ;
wire merge5_split105_bvalid ;
wire merge5_split105_bready ;


wire [IDWID-1:0] split5_merge5_arid ;
wire [31:0] split5_merge5_araddr ;
wire [7:0] split5_merge5_arlen ;
wire [EXTRAS-1:0] split5_merge5_arextras ;
wire [1:0] split5_merge5_arburst ;
wire split5_merge5_arvalid ;
wire split5_merge5_arready ;
wire [IDWID-1:0] split5_merge5_rid ;
wire [DWID-1:0] split5_merge5_rdata ;
wire [1:0] split5_merge5_rresp ;
wire split5_merge5_rlast ;
wire split5_merge5_rvalid ;
wire split5_merge5_rready ;

wire [IDWID-1:0] split5_merge5_awid ;
wire [31:0] split5_merge5_awaddr ;
wire [7:0] split5_merge5_awlen ;
wire [EXTRAS-1:0] split5_merge5_awextras ;
wire [1:0] split5_merge5_awburst ;
wire split5_merge5_awvalid ;
wire split5_merge5_awready ;
wire [DWID-1:0] split5_merge5_wdata ;
wire [WSTRB-1:0] split5_merge5_wstrb ;
wire split5_merge5_wlast ;
wire split5_merge5_wvalid ;
wire split5_merge5_wready ;
wire [IDWID-1:0] split5_merge5_bid ;
wire [1:0] split5_merge5_bresp ;
wire split5_merge5_bvalid ;
wire split5_merge5_bready ;


wire [IDWID-1:0] split6_merge5_arid ;
wire [31:0] split6_merge5_araddr ;
wire [7:0] split6_merge5_arlen ;
wire [EXTRAS-1:0] split6_merge5_arextras ;
wire [1:0] split6_merge5_arburst ;
wire split6_merge5_arvalid ;
wire split6_merge5_arready ;
wire [IDWID-1:0] split6_merge5_rid ;
wire [DWID-1:0] split6_merge5_rdata ;
wire [1:0] split6_merge5_rresp ;
wire split6_merge5_rlast ;
wire split6_merge5_rvalid ;
wire split6_merge5_rready ;

wire [IDWID-1:0] split6_merge5_awid ;
wire [31:0] split6_merge5_awaddr ;
wire [7:0] split6_merge5_awlen ;
wire [EXTRAS-1:0] split6_merge5_awextras ;
wire [1:0] split6_merge5_awburst ;
wire split6_merge5_awvalid ;
wire split6_merge5_awready ;
wire [DWID-1:0] split6_merge5_wdata ;
wire [WSTRB-1:0] split6_merge5_wstrb ;
wire split6_merge5_wlast ;
wire split6_merge5_wvalid ;
wire split6_merge5_wready ;
wire [IDWID-1:0] split6_merge5_bid ;
wire [1:0] split6_merge5_bresp ;
wire split6_merge5_bvalid ;
wire split6_merge5_bready ;


wire [IDWID-1:0] split7_merge5_arid ;
wire [31:0] split7_merge5_araddr ;
wire [7:0] split7_merge5_arlen ;
wire [EXTRAS-1:0] split7_merge5_arextras ;
wire [1:0] split7_merge5_arburst ;
wire split7_merge5_arvalid ;
wire split7_merge5_arready ;
wire [IDWID-1:0] split7_merge5_rid ;
wire [DWID-1:0] split7_merge5_rdata ;
wire [1:0] split7_merge5_rresp ;
wire split7_merge5_rlast ;
wire split7_merge5_rvalid ;
wire split7_merge5_rready ;

wire [IDWID-1:0] split7_merge5_awid ;
wire [31:0] split7_merge5_awaddr ;
wire [7:0] split7_merge5_awlen ;
wire [EXTRAS-1:0] split7_merge5_awextras ;
wire [1:0] split7_merge5_awburst ;
wire split7_merge5_awvalid ;
wire split7_merge5_awready ;
wire [DWID-1:0] split7_merge5_wdata ;
wire [WSTRB-1:0] split7_merge5_wstrb ;
wire split7_merge5_wlast ;
wire split7_merge5_wvalid ;
wire split7_merge5_wready ;
wire [IDWID-1:0] split7_merge5_bid ;
wire [1:0] split7_merge5_bresp ;
wire split7_merge5_bvalid ;
wire split7_merge5_bready ;


axi_4_merger merge5 (
     .clk(clk),.rst_n(rst_n)
    ,.araddr(merge5_split105_araddr[31:0])
    ,.arburst(merge5_split105_arburst[1:0])
    ,.arextras(merge5_split105_arextras[(EXTRAS - 1):0])
    ,.arid(merge5_split105_arid[(IDWID - 1):0])
    ,.arlen(merge5_split105_arlen[7:0])
    ,.arready(merge5_split105_arready)
    ,.arvalid(merge5_split105_arvalid)
    ,.awaddr(merge5_split105_awaddr[31:0])
    ,.awburst(merge5_split105_awburst[1:0])
    ,.awextras(merge5_split105_awextras[(EXTRAS - 1):0])
    ,.awid(merge5_split105_awid[3:0])
    ,.awlen(merge5_split105_awlen[7:0])
    ,.awready(merge5_split105_awready)
    ,.awvalid(merge5_split105_awvalid)
    ,.bid(merge5_split105_bid[(IDWID - 1):0])
    ,.bready(merge5_split105_bready)
    ,.bresp(merge5_split105_bresp[1:0])
    ,.bvalid(merge5_split105_bvalid)
    ,.rid(merge5_split105_rid[(IDWID - 1):0])
    ,.rlast(merge5_split105_rlast)
    ,.rready(merge5_split105_rready)
    ,.rresp(merge5_split105_rresp[1:0])
    ,.rvalid(merge5_split105_rvalid)
    ,.rdata(merge5_split105_rdata[(DWID - 1):0])
    ,.wdata(merge5_split105_wdata[(DWID - 1):0])
    ,.wlast(merge5_split105_wlast)
    ,.wready(merge5_split105_wready)
    ,.wstrb(merge5_split105_wstrb[(WSTRB - 1):0])
    ,.wvalid(merge5_split105_wvalid)


    ,.a_araddr(split4_merge5_araddr[31:0])
    ,.a_arburst(split4_merge5_arburst[1:0])
    ,.a_arextras(split4_merge5_arextras[(EXTRAS - 1):0])
    ,.a_arid(split4_merge5_arid[(IDWID - 1):0])
    ,.a_arlen(split4_merge5_arlen[7:0])
    ,.a_arready(split4_merge5_arready)
    ,.a_arvalid(split4_merge5_arvalid)
    ,.a_awaddr(split4_merge5_awaddr[31:0])
    ,.a_awburst(split4_merge5_awburst[1:0])
    ,.a_awextras(split4_merge5_awextras[(EXTRAS - 1):0])
    ,.a_awid(split4_merge5_awid[(IDWID - 1):0])
    ,.a_awlen(split4_merge5_awlen[7:0])
    ,.a_awready(split4_merge5_awready)
    ,.a_awvalid(split4_merge5_awvalid)
    ,.a_bid(split4_merge5_bid[(IDWID - 1):0])
    ,.a_bready(split4_merge5_bready)
    ,.a_bresp(split4_merge5_bresp[1:0])
    ,.a_bvalid(split4_merge5_bvalid)
    ,.a_rdata(split4_merge5_rdata[(DWID - 1):0])
    ,.a_rid(split4_merge5_rid[(IDWID - 1):0])
    ,.a_rlast(split4_merge5_rlast)
    ,.a_rready(split4_merge5_rready)
    ,.a_rresp(split4_merge5_rresp[1:0])
    ,.a_rvalid(split4_merge5_rvalid)
    ,.a_wdata(split4_merge5_wdata[(DWID - 1):0])
    ,.a_wlast(split4_merge5_wlast)
    ,.a_wready(split4_merge5_wready)
    ,.a_wstrb(split4_merge5_wstrb[(WSTRB - 1):0])
    ,.a_wvalid(split4_merge5_wvalid)

    ,.b_araddr(split5_merge5_araddr[31:0])
    ,.b_arburst(split5_merge5_arburst[1:0])
    ,.b_arextras(split5_merge5_arextras[(EXTRAS - 1):0])
    ,.b_arid(split5_merge5_arid[(IDWID - 1):0])
    ,.b_arlen(split5_merge5_arlen[7:0])
    ,.b_arready(split5_merge5_arready)
    ,.b_arvalid(split5_merge5_arvalid)
    ,.b_awaddr(split5_merge5_awaddr[31:0])
    ,.b_awburst(split5_merge5_awburst[1:0])
    ,.b_awextras(split5_merge5_awextras[(EXTRAS - 1):0])
    ,.b_awid(split5_merge5_awid[(IDWID - 1):0])
    ,.b_awlen(split5_merge5_awlen[7:0])
    ,.b_awready(split5_merge5_awready)
    ,.b_awvalid(split5_merge5_awvalid)
    ,.b_bid(split5_merge5_bid[(IDWID - 1):0])
    ,.b_bready(split5_merge5_bready)
    ,.b_bresp(split5_merge5_bresp[1:0])
    ,.b_bvalid(split5_merge5_bvalid)
    ,.b_rdata(split5_merge5_rdata[(DWID - 1):0])
    ,.b_rid(split5_merge5_rid[(IDWID - 1):0])
    ,.b_rlast(split5_merge5_rlast)
    ,.b_rready(split5_merge5_rready)
    ,.b_rresp(split5_merge5_rresp[1:0])
    ,.b_rvalid(split5_merge5_rvalid)
    ,.b_wdata(split5_merge5_wdata[(DWID - 1):0])
    ,.b_wlast(split5_merge5_wlast)
    ,.b_wready(split5_merge5_wready)
    ,.b_wstrb(split5_merge5_wstrb[(WSTRB - 1):0])
    ,.b_wvalid(split5_merge5_wvalid)

    ,.c_araddr(split6_merge5_araddr[31:0])
    ,.c_arburst(split6_merge5_arburst[1:0])
    ,.c_arextras(split6_merge5_arextras[(EXTRAS - 1):0])
    ,.c_arid(split6_merge5_arid[(IDWID - 1):0])
    ,.c_arlen(split6_merge5_arlen[7:0])
    ,.c_arready(split6_merge5_arready)
    ,.c_arvalid(split6_merge5_arvalid)
    ,.c_awaddr(split6_merge5_awaddr[31:0])
    ,.c_awburst(split6_merge5_awburst[1:0])
    ,.c_awextras(split6_merge5_awextras[(EXTRAS - 1):0])
    ,.c_awid(split6_merge5_awid[(IDWID - 1):0])
    ,.c_awlen(split6_merge5_awlen[7:0])
    ,.c_awready(split6_merge5_awready)
    ,.c_awvalid(split6_merge5_awvalid)
    ,.c_bid(split6_merge5_bid[(IDWID - 1):0])
    ,.c_bready(split6_merge5_bready)
    ,.c_bresp(split6_merge5_bresp[1:0])
    ,.c_bvalid(split6_merge5_bvalid)
    ,.c_rdata(split6_merge5_rdata[(DWID - 1):0])
    ,.c_rid(split6_merge5_rid[(IDWID - 1):0])
    ,.c_rlast(split6_merge5_rlast)
    ,.c_rready(split6_merge5_rready)
    ,.c_rresp(split6_merge5_rresp[1:0])
    ,.c_rvalid(split6_merge5_rvalid)
    ,.c_wdata(split6_merge5_wdata[(DWID - 1):0])
    ,.c_wlast(split6_merge5_wlast)
    ,.c_wready(split6_merge5_wready)
    ,.c_wstrb(split6_merge5_wstrb[(WSTRB - 1):0])
    ,.c_wvalid(split6_merge5_wvalid)

    ,.d_araddr(split7_merge5_araddr[31:0])
    ,.d_arburst(split7_merge5_arburst[1:0])
    ,.d_arextras(split7_merge5_arextras[(EXTRAS - 1):0])
    ,.d_arid(split7_merge5_arid[(IDWID - 1):0])
    ,.d_arlen(split7_merge5_arlen[7:0])
    ,.d_arready(split7_merge5_arready)
    ,.d_arvalid(split7_merge5_arvalid)
    ,.d_awaddr(split7_merge5_awaddr[31:0])
    ,.d_awburst(split7_merge5_awburst[1:0])
    ,.d_awextras(split7_merge5_awextras[(EXTRAS - 1):0])
    ,.d_awid(split7_merge5_awid[(IDWID - 1):0])
    ,.d_awlen(split7_merge5_awlen[7:0])
    ,.d_awready(split7_merge5_awready)
    ,.d_awvalid(split7_merge5_awvalid)
    ,.d_bid(split7_merge5_bid[(IDWID - 1):0])
    ,.d_bready(split7_merge5_bready)
    ,.d_bresp(split7_merge5_bresp[1:0])
    ,.d_bvalid(split7_merge5_bvalid)
    ,.d_rdata(split7_merge5_rdata[(DWID - 1):0])
    ,.d_rid(split7_merge5_rid[(IDWID - 1):0])
    ,.d_rlast(split7_merge5_rlast)
    ,.d_rready(split7_merge5_rready)
    ,.d_rresp(split7_merge5_rresp[1:0])
    ,.d_rvalid(split7_merge5_rvalid)
    ,.d_wdata(split7_merge5_wdata[(DWID - 1):0])
    ,.d_wlast(split7_merge5_wlast)
    ,.d_wready(split7_merge5_wready)
    ,.d_wstrb(split7_merge5_wstrb[(WSTRB - 1):0])
    ,.d_wvalid(split7_merge5_wvalid)
);


wire [IDWID-1:0] merge6_split106_arid ;
wire [31:0] merge6_split106_araddr ;
wire [7:0] merge6_split106_arlen ;
wire [EXTRAS-1:0] merge6_split106_arextras ;
wire [1:0] merge6_split106_arburst ;
wire merge6_split106_arvalid ;
wire merge6_split106_arready ;
wire [IDWID-1:0] merge6_split106_rid ;
wire [DWID-1:0] merge6_split106_rdata ;
wire [1:0] merge6_split106_rresp ;
wire merge6_split106_rlast ;
wire merge6_split106_rvalid ;
wire merge6_split106_rready ;

wire [IDWID-1:0] merge6_split106_awid ;
wire [31:0] merge6_split106_awaddr ;
wire [7:0] merge6_split106_awlen ;
wire [EXTRAS-1:0] merge6_split106_awextras ;
wire [1:0] merge6_split106_awburst ;
wire merge6_split106_awvalid ;
wire merge6_split106_awready ;
wire [DWID-1:0] merge6_split106_wdata ;
wire [WSTRB-1:0] merge6_split106_wstrb ;
wire merge6_split106_wlast ;
wire merge6_split106_wvalid ;
wire merge6_split106_wready ;
wire [IDWID-1:0] merge6_split106_bid ;
wire [1:0] merge6_split106_bresp ;
wire merge6_split106_bvalid ;
wire merge6_split106_bready ;


wire [IDWID-1:0] split5_merge6_arid ;
wire [31:0] split5_merge6_araddr ;
wire [7:0] split5_merge6_arlen ;
wire [EXTRAS-1:0] split5_merge6_arextras ;
wire [1:0] split5_merge6_arburst ;
wire split5_merge6_arvalid ;
wire split5_merge6_arready ;
wire [IDWID-1:0] split5_merge6_rid ;
wire [DWID-1:0] split5_merge6_rdata ;
wire [1:0] split5_merge6_rresp ;
wire split5_merge6_rlast ;
wire split5_merge6_rvalid ;
wire split5_merge6_rready ;

wire [IDWID-1:0] split5_merge6_awid ;
wire [31:0] split5_merge6_awaddr ;
wire [7:0] split5_merge6_awlen ;
wire [EXTRAS-1:0] split5_merge6_awextras ;
wire [1:0] split5_merge6_awburst ;
wire split5_merge6_awvalid ;
wire split5_merge6_awready ;
wire [DWID-1:0] split5_merge6_wdata ;
wire [WSTRB-1:0] split5_merge6_wstrb ;
wire split5_merge6_wlast ;
wire split5_merge6_wvalid ;
wire split5_merge6_wready ;
wire [IDWID-1:0] split5_merge6_bid ;
wire [1:0] split5_merge6_bresp ;
wire split5_merge6_bvalid ;
wire split5_merge6_bready ;


wire [IDWID-1:0] split6_merge6_arid ;
wire [31:0] split6_merge6_araddr ;
wire [7:0] split6_merge6_arlen ;
wire [EXTRAS-1:0] split6_merge6_arextras ;
wire [1:0] split6_merge6_arburst ;
wire split6_merge6_arvalid ;
wire split6_merge6_arready ;
wire [IDWID-1:0] split6_merge6_rid ;
wire [DWID-1:0] split6_merge6_rdata ;
wire [1:0] split6_merge6_rresp ;
wire split6_merge6_rlast ;
wire split6_merge6_rvalid ;
wire split6_merge6_rready ;

wire [IDWID-1:0] split6_merge6_awid ;
wire [31:0] split6_merge6_awaddr ;
wire [7:0] split6_merge6_awlen ;
wire [EXTRAS-1:0] split6_merge6_awextras ;
wire [1:0] split6_merge6_awburst ;
wire split6_merge6_awvalid ;
wire split6_merge6_awready ;
wire [DWID-1:0] split6_merge6_wdata ;
wire [WSTRB-1:0] split6_merge6_wstrb ;
wire split6_merge6_wlast ;
wire split6_merge6_wvalid ;
wire split6_merge6_wready ;
wire [IDWID-1:0] split6_merge6_bid ;
wire [1:0] split6_merge6_bresp ;
wire split6_merge6_bvalid ;
wire split6_merge6_bready ;


wire [IDWID-1:0] split7_merge6_arid ;
wire [31:0] split7_merge6_araddr ;
wire [7:0] split7_merge6_arlen ;
wire [EXTRAS-1:0] split7_merge6_arextras ;
wire [1:0] split7_merge6_arburst ;
wire split7_merge6_arvalid ;
wire split7_merge6_arready ;
wire [IDWID-1:0] split7_merge6_rid ;
wire [DWID-1:0] split7_merge6_rdata ;
wire [1:0] split7_merge6_rresp ;
wire split7_merge6_rlast ;
wire split7_merge6_rvalid ;
wire split7_merge6_rready ;

wire [IDWID-1:0] split7_merge6_awid ;
wire [31:0] split7_merge6_awaddr ;
wire [7:0] split7_merge6_awlen ;
wire [EXTRAS-1:0] split7_merge6_awextras ;
wire [1:0] split7_merge6_awburst ;
wire split7_merge6_awvalid ;
wire split7_merge6_awready ;
wire [DWID-1:0] split7_merge6_wdata ;
wire [WSTRB-1:0] split7_merge6_wstrb ;
wire split7_merge6_wlast ;
wire split7_merge6_wvalid ;
wire split7_merge6_wready ;
wire [IDWID-1:0] split7_merge6_bid ;
wire [1:0] split7_merge6_bresp ;
wire split7_merge6_bvalid ;
wire split7_merge6_bready ;


axi_4_merger merge6 (
     .clk(clk),.rst_n(rst_n)
    ,.araddr(merge6_split106_araddr[31:0])
    ,.arburst(merge6_split106_arburst[1:0])
    ,.arextras(merge6_split106_arextras[(EXTRAS - 1):0])
    ,.arid(merge6_split106_arid[(IDWID - 1):0])
    ,.arlen(merge6_split106_arlen[7:0])
    ,.arready(merge6_split106_arready)
    ,.arvalid(merge6_split106_arvalid)
    ,.awaddr(merge6_split106_awaddr[31:0])
    ,.awburst(merge6_split106_awburst[1:0])
    ,.awextras(merge6_split106_awextras[(EXTRAS - 1):0])
    ,.awid(merge6_split106_awid[3:0])
    ,.awlen(merge6_split106_awlen[7:0])
    ,.awready(merge6_split106_awready)
    ,.awvalid(merge6_split106_awvalid)
    ,.bid(merge6_split106_bid[(IDWID - 1):0])
    ,.bready(merge6_split106_bready)
    ,.bresp(merge6_split106_bresp[1:0])
    ,.bvalid(merge6_split106_bvalid)
    ,.rid(merge6_split106_rid[(IDWID - 1):0])
    ,.rlast(merge6_split106_rlast)
    ,.rready(merge6_split106_rready)
    ,.rresp(merge6_split106_rresp[1:0])
    ,.rvalid(merge6_split106_rvalid)
    ,.rdata(merge6_split106_rdata[(DWID - 1):0])
    ,.wdata(merge6_split106_wdata[(DWID - 1):0])
    ,.wlast(merge6_split106_wlast)
    ,.wready(merge6_split106_wready)
    ,.wstrb(merge6_split106_wstrb[(WSTRB - 1):0])
    ,.wvalid(merge6_split106_wvalid)


    ,.a_araddr(split4_merge6_araddr[31:0])
    ,.a_arburst(split4_merge6_arburst[1:0])
    ,.a_arextras(split4_merge6_arextras[(EXTRAS - 1):0])
    ,.a_arid(split4_merge6_arid[(IDWID - 1):0])
    ,.a_arlen(split4_merge6_arlen[7:0])
    ,.a_arready(split4_merge6_arready)
    ,.a_arvalid(split4_merge6_arvalid)
    ,.a_awaddr(split4_merge6_awaddr[31:0])
    ,.a_awburst(split4_merge6_awburst[1:0])
    ,.a_awextras(split4_merge6_awextras[(EXTRAS - 1):0])
    ,.a_awid(split4_merge6_awid[(IDWID - 1):0])
    ,.a_awlen(split4_merge6_awlen[7:0])
    ,.a_awready(split4_merge6_awready)
    ,.a_awvalid(split4_merge6_awvalid)
    ,.a_bid(split4_merge6_bid[(IDWID - 1):0])
    ,.a_bready(split4_merge6_bready)
    ,.a_bresp(split4_merge6_bresp[1:0])
    ,.a_bvalid(split4_merge6_bvalid)
    ,.a_rdata(split4_merge6_rdata[(DWID - 1):0])
    ,.a_rid(split4_merge6_rid[(IDWID - 1):0])
    ,.a_rlast(split4_merge6_rlast)
    ,.a_rready(split4_merge6_rready)
    ,.a_rresp(split4_merge6_rresp[1:0])
    ,.a_rvalid(split4_merge6_rvalid)
    ,.a_wdata(split4_merge6_wdata[(DWID - 1):0])
    ,.a_wlast(split4_merge6_wlast)
    ,.a_wready(split4_merge6_wready)
    ,.a_wstrb(split4_merge6_wstrb[(WSTRB - 1):0])
    ,.a_wvalid(split4_merge6_wvalid)

    ,.b_araddr(split5_merge6_araddr[31:0])
    ,.b_arburst(split5_merge6_arburst[1:0])
    ,.b_arextras(split5_merge6_arextras[(EXTRAS - 1):0])
    ,.b_arid(split5_merge6_arid[(IDWID - 1):0])
    ,.b_arlen(split5_merge6_arlen[7:0])
    ,.b_arready(split5_merge6_arready)
    ,.b_arvalid(split5_merge6_arvalid)
    ,.b_awaddr(split5_merge6_awaddr[31:0])
    ,.b_awburst(split5_merge6_awburst[1:0])
    ,.b_awextras(split5_merge6_awextras[(EXTRAS - 1):0])
    ,.b_awid(split5_merge6_awid[(IDWID - 1):0])
    ,.b_awlen(split5_merge6_awlen[7:0])
    ,.b_awready(split5_merge6_awready)
    ,.b_awvalid(split5_merge6_awvalid)
    ,.b_bid(split5_merge6_bid[(IDWID - 1):0])
    ,.b_bready(split5_merge6_bready)
    ,.b_bresp(split5_merge6_bresp[1:0])
    ,.b_bvalid(split5_merge6_bvalid)
    ,.b_rdata(split5_merge6_rdata[(DWID - 1):0])
    ,.b_rid(split5_merge6_rid[(IDWID - 1):0])
    ,.b_rlast(split5_merge6_rlast)
    ,.b_rready(split5_merge6_rready)
    ,.b_rresp(split5_merge6_rresp[1:0])
    ,.b_rvalid(split5_merge6_rvalid)
    ,.b_wdata(split5_merge6_wdata[(DWID - 1):0])
    ,.b_wlast(split5_merge6_wlast)
    ,.b_wready(split5_merge6_wready)
    ,.b_wstrb(split5_merge6_wstrb[(WSTRB - 1):0])
    ,.b_wvalid(split5_merge6_wvalid)

    ,.c_araddr(split6_merge6_araddr[31:0])
    ,.c_arburst(split6_merge6_arburst[1:0])
    ,.c_arextras(split6_merge6_arextras[(EXTRAS - 1):0])
    ,.c_arid(split6_merge6_arid[(IDWID - 1):0])
    ,.c_arlen(split6_merge6_arlen[7:0])
    ,.c_arready(split6_merge6_arready)
    ,.c_arvalid(split6_merge6_arvalid)
    ,.c_awaddr(split6_merge6_awaddr[31:0])
    ,.c_awburst(split6_merge6_awburst[1:0])
    ,.c_awextras(split6_merge6_awextras[(EXTRAS - 1):0])
    ,.c_awid(split6_merge6_awid[(IDWID - 1):0])
    ,.c_awlen(split6_merge6_awlen[7:0])
    ,.c_awready(split6_merge6_awready)
    ,.c_awvalid(split6_merge6_awvalid)
    ,.c_bid(split6_merge6_bid[(IDWID - 1):0])
    ,.c_bready(split6_merge6_bready)
    ,.c_bresp(split6_merge6_bresp[1:0])
    ,.c_bvalid(split6_merge6_bvalid)
    ,.c_rdata(split6_merge6_rdata[(DWID - 1):0])
    ,.c_rid(split6_merge6_rid[(IDWID - 1):0])
    ,.c_rlast(split6_merge6_rlast)
    ,.c_rready(split6_merge6_rready)
    ,.c_rresp(split6_merge6_rresp[1:0])
    ,.c_rvalid(split6_merge6_rvalid)
    ,.c_wdata(split6_merge6_wdata[(DWID - 1):0])
    ,.c_wlast(split6_merge6_wlast)
    ,.c_wready(split6_merge6_wready)
    ,.c_wstrb(split6_merge6_wstrb[(WSTRB - 1):0])
    ,.c_wvalid(split6_merge6_wvalid)

    ,.d_araddr(split7_merge6_araddr[31:0])
    ,.d_arburst(split7_merge6_arburst[1:0])
    ,.d_arextras(split7_merge6_arextras[(EXTRAS - 1):0])
    ,.d_arid(split7_merge6_arid[(IDWID - 1):0])
    ,.d_arlen(split7_merge6_arlen[7:0])
    ,.d_arready(split7_merge6_arready)
    ,.d_arvalid(split7_merge6_arvalid)
    ,.d_awaddr(split7_merge6_awaddr[31:0])
    ,.d_awburst(split7_merge6_awburst[1:0])
    ,.d_awextras(split7_merge6_awextras[(EXTRAS - 1):0])
    ,.d_awid(split7_merge6_awid[(IDWID - 1):0])
    ,.d_awlen(split7_merge6_awlen[7:0])
    ,.d_awready(split7_merge6_awready)
    ,.d_awvalid(split7_merge6_awvalid)
    ,.d_bid(split7_merge6_bid[(IDWID - 1):0])
    ,.d_bready(split7_merge6_bready)
    ,.d_bresp(split7_merge6_bresp[1:0])
    ,.d_bvalid(split7_merge6_bvalid)
    ,.d_rdata(split7_merge6_rdata[(DWID - 1):0])
    ,.d_rid(split7_merge6_rid[(IDWID - 1):0])
    ,.d_rlast(split7_merge6_rlast)
    ,.d_rready(split7_merge6_rready)
    ,.d_rresp(split7_merge6_rresp[1:0])
    ,.d_rvalid(split7_merge6_rvalid)
    ,.d_wdata(split7_merge6_wdata[(DWID - 1):0])
    ,.d_wlast(split7_merge6_wlast)
    ,.d_wready(split7_merge6_wready)
    ,.d_wstrb(split7_merge6_wstrb[(WSTRB - 1):0])
    ,.d_wvalid(split7_merge6_wvalid)
);


wire [IDWID-1:0] merge7_split107_arid ;
wire [31:0] merge7_split107_araddr ;
wire [7:0] merge7_split107_arlen ;
wire [EXTRAS-1:0] merge7_split107_arextras ;
wire [1:0] merge7_split107_arburst ;
wire merge7_split107_arvalid ;
wire merge7_split107_arready ;
wire [IDWID-1:0] merge7_split107_rid ;
wire [DWID-1:0] merge7_split107_rdata ;
wire [1:0] merge7_split107_rresp ;
wire merge7_split107_rlast ;
wire merge7_split107_rvalid ;
wire merge7_split107_rready ;

wire [IDWID-1:0] merge7_split107_awid ;
wire [31:0] merge7_split107_awaddr ;
wire [7:0] merge7_split107_awlen ;
wire [EXTRAS-1:0] merge7_split107_awextras ;
wire [1:0] merge7_split107_awburst ;
wire merge7_split107_awvalid ;
wire merge7_split107_awready ;
wire [DWID-1:0] merge7_split107_wdata ;
wire [WSTRB-1:0] merge7_split107_wstrb ;
wire merge7_split107_wlast ;
wire merge7_split107_wvalid ;
wire merge7_split107_wready ;
wire [IDWID-1:0] merge7_split107_bid ;
wire [1:0] merge7_split107_bresp ;
wire merge7_split107_bvalid ;
wire merge7_split107_bready ;


wire [IDWID-1:0] split5_merge7_arid ;
wire [31:0] split5_merge7_araddr ;
wire [7:0] split5_merge7_arlen ;
wire [EXTRAS-1:0] split5_merge7_arextras ;
wire [1:0] split5_merge7_arburst ;
wire split5_merge7_arvalid ;
wire split5_merge7_arready ;
wire [IDWID-1:0] split5_merge7_rid ;
wire [DWID-1:0] split5_merge7_rdata ;
wire [1:0] split5_merge7_rresp ;
wire split5_merge7_rlast ;
wire split5_merge7_rvalid ;
wire split5_merge7_rready ;

wire [IDWID-1:0] split5_merge7_awid ;
wire [31:0] split5_merge7_awaddr ;
wire [7:0] split5_merge7_awlen ;
wire [EXTRAS-1:0] split5_merge7_awextras ;
wire [1:0] split5_merge7_awburst ;
wire split5_merge7_awvalid ;
wire split5_merge7_awready ;
wire [DWID-1:0] split5_merge7_wdata ;
wire [WSTRB-1:0] split5_merge7_wstrb ;
wire split5_merge7_wlast ;
wire split5_merge7_wvalid ;
wire split5_merge7_wready ;
wire [IDWID-1:0] split5_merge7_bid ;
wire [1:0] split5_merge7_bresp ;
wire split5_merge7_bvalid ;
wire split5_merge7_bready ;


wire [IDWID-1:0] split6_merge7_arid ;
wire [31:0] split6_merge7_araddr ;
wire [7:0] split6_merge7_arlen ;
wire [EXTRAS-1:0] split6_merge7_arextras ;
wire [1:0] split6_merge7_arburst ;
wire split6_merge7_arvalid ;
wire split6_merge7_arready ;
wire [IDWID-1:0] split6_merge7_rid ;
wire [DWID-1:0] split6_merge7_rdata ;
wire [1:0] split6_merge7_rresp ;
wire split6_merge7_rlast ;
wire split6_merge7_rvalid ;
wire split6_merge7_rready ;

wire [IDWID-1:0] split6_merge7_awid ;
wire [31:0] split6_merge7_awaddr ;
wire [7:0] split6_merge7_awlen ;
wire [EXTRAS-1:0] split6_merge7_awextras ;
wire [1:0] split6_merge7_awburst ;
wire split6_merge7_awvalid ;
wire split6_merge7_awready ;
wire [DWID-1:0] split6_merge7_wdata ;
wire [WSTRB-1:0] split6_merge7_wstrb ;
wire split6_merge7_wlast ;
wire split6_merge7_wvalid ;
wire split6_merge7_wready ;
wire [IDWID-1:0] split6_merge7_bid ;
wire [1:0] split6_merge7_bresp ;
wire split6_merge7_bvalid ;
wire split6_merge7_bready ;


wire [IDWID-1:0] split7_merge7_arid ;
wire [31:0] split7_merge7_araddr ;
wire [7:0] split7_merge7_arlen ;
wire [EXTRAS-1:0] split7_merge7_arextras ;
wire [1:0] split7_merge7_arburst ;
wire split7_merge7_arvalid ;
wire split7_merge7_arready ;
wire [IDWID-1:0] split7_merge7_rid ;
wire [DWID-1:0] split7_merge7_rdata ;
wire [1:0] split7_merge7_rresp ;
wire split7_merge7_rlast ;
wire split7_merge7_rvalid ;
wire split7_merge7_rready ;

wire [IDWID-1:0] split7_merge7_awid ;
wire [31:0] split7_merge7_awaddr ;
wire [7:0] split7_merge7_awlen ;
wire [EXTRAS-1:0] split7_merge7_awextras ;
wire [1:0] split7_merge7_awburst ;
wire split7_merge7_awvalid ;
wire split7_merge7_awready ;
wire [DWID-1:0] split7_merge7_wdata ;
wire [WSTRB-1:0] split7_merge7_wstrb ;
wire split7_merge7_wlast ;
wire split7_merge7_wvalid ;
wire split7_merge7_wready ;
wire [IDWID-1:0] split7_merge7_bid ;
wire [1:0] split7_merge7_bresp ;
wire split7_merge7_bvalid ;
wire split7_merge7_bready ;


axi_4_merger merge7 (
     .clk(clk),.rst_n(rst_n)
    ,.araddr(merge7_split107_araddr[31:0])
    ,.arburst(merge7_split107_arburst[1:0])
    ,.arextras(merge7_split107_arextras[(EXTRAS - 1):0])
    ,.arid(merge7_split107_arid[(IDWID - 1):0])
    ,.arlen(merge7_split107_arlen[7:0])
    ,.arready(merge7_split107_arready)
    ,.arvalid(merge7_split107_arvalid)
    ,.awaddr(merge7_split107_awaddr[31:0])
    ,.awburst(merge7_split107_awburst[1:0])
    ,.awextras(merge7_split107_awextras[(EXTRAS - 1):0])
    ,.awid(merge7_split107_awid[3:0])
    ,.awlen(merge7_split107_awlen[7:0])
    ,.awready(merge7_split107_awready)
    ,.awvalid(merge7_split107_awvalid)
    ,.bid(merge7_split107_bid[(IDWID - 1):0])
    ,.bready(merge7_split107_bready)
    ,.bresp(merge7_split107_bresp[1:0])
    ,.bvalid(merge7_split107_bvalid)
    ,.rid(merge7_split107_rid[(IDWID - 1):0])
    ,.rlast(merge7_split107_rlast)
    ,.rready(merge7_split107_rready)
    ,.rresp(merge7_split107_rresp[1:0])
    ,.rvalid(merge7_split107_rvalid)
    ,.rdata(merge7_split107_rdata[(DWID - 1):0])
    ,.wdata(merge7_split107_wdata[(DWID - 1):0])
    ,.wlast(merge7_split107_wlast)
    ,.wready(merge7_split107_wready)
    ,.wstrb(merge7_split107_wstrb[(WSTRB - 1):0])
    ,.wvalid(merge7_split107_wvalid)


    ,.a_araddr(split4_merge7_araddr[31:0])
    ,.a_arburst(split4_merge7_arburst[1:0])
    ,.a_arextras(split4_merge7_arextras[(EXTRAS - 1):0])
    ,.a_arid(split4_merge7_arid[(IDWID - 1):0])
    ,.a_arlen(split4_merge7_arlen[7:0])
    ,.a_arready(split4_merge7_arready)
    ,.a_arvalid(split4_merge7_arvalid)
    ,.a_awaddr(split4_merge7_awaddr[31:0])
    ,.a_awburst(split4_merge7_awburst[1:0])
    ,.a_awextras(split4_merge7_awextras[(EXTRAS - 1):0])
    ,.a_awid(split4_merge7_awid[(IDWID - 1):0])
    ,.a_awlen(split4_merge7_awlen[7:0])
    ,.a_awready(split4_merge7_awready)
    ,.a_awvalid(split4_merge7_awvalid)
    ,.a_bid(split4_merge7_bid[(IDWID - 1):0])
    ,.a_bready(split4_merge7_bready)
    ,.a_bresp(split4_merge7_bresp[1:0])
    ,.a_bvalid(split4_merge7_bvalid)
    ,.a_rdata(split4_merge7_rdata[(DWID - 1):0])
    ,.a_rid(split4_merge7_rid[(IDWID - 1):0])
    ,.a_rlast(split4_merge7_rlast)
    ,.a_rready(split4_merge7_rready)
    ,.a_rresp(split4_merge7_rresp[1:0])
    ,.a_rvalid(split4_merge7_rvalid)
    ,.a_wdata(split4_merge7_wdata[(DWID - 1):0])
    ,.a_wlast(split4_merge7_wlast)
    ,.a_wready(split4_merge7_wready)
    ,.a_wstrb(split4_merge7_wstrb[(WSTRB - 1):0])
    ,.a_wvalid(split4_merge7_wvalid)

    ,.b_araddr(split5_merge7_araddr[31:0])
    ,.b_arburst(split5_merge7_arburst[1:0])
    ,.b_arextras(split5_merge7_arextras[(EXTRAS - 1):0])
    ,.b_arid(split5_merge7_arid[(IDWID - 1):0])
    ,.b_arlen(split5_merge7_arlen[7:0])
    ,.b_arready(split5_merge7_arready)
    ,.b_arvalid(split5_merge7_arvalid)
    ,.b_awaddr(split5_merge7_awaddr[31:0])
    ,.b_awburst(split5_merge7_awburst[1:0])
    ,.b_awextras(split5_merge7_awextras[(EXTRAS - 1):0])
    ,.b_awid(split5_merge7_awid[(IDWID - 1):0])
    ,.b_awlen(split5_merge7_awlen[7:0])
    ,.b_awready(split5_merge7_awready)
    ,.b_awvalid(split5_merge7_awvalid)
    ,.b_bid(split5_merge7_bid[(IDWID - 1):0])
    ,.b_bready(split5_merge7_bready)
    ,.b_bresp(split5_merge7_bresp[1:0])
    ,.b_bvalid(split5_merge7_bvalid)
    ,.b_rdata(split5_merge7_rdata[(DWID - 1):0])
    ,.b_rid(split5_merge7_rid[(IDWID - 1):0])
    ,.b_rlast(split5_merge7_rlast)
    ,.b_rready(split5_merge7_rready)
    ,.b_rresp(split5_merge7_rresp[1:0])
    ,.b_rvalid(split5_merge7_rvalid)
    ,.b_wdata(split5_merge7_wdata[(DWID - 1):0])
    ,.b_wlast(split5_merge7_wlast)
    ,.b_wready(split5_merge7_wready)
    ,.b_wstrb(split5_merge7_wstrb[(WSTRB - 1):0])
    ,.b_wvalid(split5_merge7_wvalid)

    ,.c_araddr(split6_merge7_araddr[31:0])
    ,.c_arburst(split6_merge7_arburst[1:0])
    ,.c_arextras(split6_merge7_arextras[(EXTRAS - 1):0])
    ,.c_arid(split6_merge7_arid[(IDWID - 1):0])
    ,.c_arlen(split6_merge7_arlen[7:0])
    ,.c_arready(split6_merge7_arready)
    ,.c_arvalid(split6_merge7_arvalid)
    ,.c_awaddr(split6_merge7_awaddr[31:0])
    ,.c_awburst(split6_merge7_awburst[1:0])
    ,.c_awextras(split6_merge7_awextras[(EXTRAS - 1):0])
    ,.c_awid(split6_merge7_awid[(IDWID - 1):0])
    ,.c_awlen(split6_merge7_awlen[7:0])
    ,.c_awready(split6_merge7_awready)
    ,.c_awvalid(split6_merge7_awvalid)
    ,.c_bid(split6_merge7_bid[(IDWID - 1):0])
    ,.c_bready(split6_merge7_bready)
    ,.c_bresp(split6_merge7_bresp[1:0])
    ,.c_bvalid(split6_merge7_bvalid)
    ,.c_rdata(split6_merge7_rdata[(DWID - 1):0])
    ,.c_rid(split6_merge7_rid[(IDWID - 1):0])
    ,.c_rlast(split6_merge7_rlast)
    ,.c_rready(split6_merge7_rready)
    ,.c_rresp(split6_merge7_rresp[1:0])
    ,.c_rvalid(split6_merge7_rvalid)
    ,.c_wdata(split6_merge7_wdata[(DWID - 1):0])
    ,.c_wlast(split6_merge7_wlast)
    ,.c_wready(split6_merge7_wready)
    ,.c_wstrb(split6_merge7_wstrb[(WSTRB - 1):0])
    ,.c_wvalid(split6_merge7_wvalid)

    ,.d_araddr(split7_merge7_araddr[31:0])
    ,.d_arburst(split7_merge7_arburst[1:0])
    ,.d_arextras(split7_merge7_arextras[(EXTRAS - 1):0])
    ,.d_arid(split7_merge7_arid[(IDWID - 1):0])
    ,.d_arlen(split7_merge7_arlen[7:0])
    ,.d_arready(split7_merge7_arready)
    ,.d_arvalid(split7_merge7_arvalid)
    ,.d_awaddr(split7_merge7_awaddr[31:0])
    ,.d_awburst(split7_merge7_awburst[1:0])
    ,.d_awextras(split7_merge7_awextras[(EXTRAS - 1):0])
    ,.d_awid(split7_merge7_awid[(IDWID - 1):0])
    ,.d_awlen(split7_merge7_awlen[7:0])
    ,.d_awready(split7_merge7_awready)
    ,.d_awvalid(split7_merge7_awvalid)
    ,.d_bid(split7_merge7_bid[(IDWID - 1):0])
    ,.d_bready(split7_merge7_bready)
    ,.d_bresp(split7_merge7_bresp[1:0])
    ,.d_bvalid(split7_merge7_bvalid)
    ,.d_rdata(split7_merge7_rdata[(DWID - 1):0])
    ,.d_rid(split7_merge7_rid[(IDWID - 1):0])
    ,.d_rlast(split7_merge7_rlast)
    ,.d_rready(split7_merge7_rready)
    ,.d_rresp(split7_merge7_rresp[1:0])
    ,.d_rvalid(split7_merge7_rvalid)
    ,.d_wdata(split7_merge7_wdata[(DWID - 1):0])
    ,.d_wlast(split7_merge7_wlast)
    ,.d_wready(split7_merge7_wready)
    ,.d_wstrb(split7_merge7_wstrb[(WSTRB - 1):0])
    ,.d_wvalid(split7_merge7_wvalid)
);


axi_4_splitter split5 (
     .clk(clk) ,.rst_n(rst_n)

    ,.araddr(mst5_araddr[31:0])
    ,.arburst(mst5_arburst[1:0])
    ,.arextras(mst5_arextras[(EXTRAS - 1):0])
    ,.arid(mst5_arid[(IDWID - 1):0])
    ,.arlen(mst5_arlen[7:0])
    ,.arready(mst5_arready)
    ,.arvalid(mst5_arvalid)
    ,.awaddr(mst5_awaddr[31:0])
    ,.awburst(mst5_awburst[1:0])
    ,.awextras(mst5_awextras[(EXTRAS - 1):0])
    ,.awid(mst5_awid[3:0])
    ,.awlen(mst5_awlen[7:0])
    ,.awready(mst5_awready)
    ,.awvalid(mst5_awvalid)
    ,.bid(mst5_bid[(IDWID - 1):0])
    ,.bready(mst5_bready)
    ,.bresp(mst5_bresp[1:0])
    ,.bvalid(mst5_bvalid)
    ,.rdata(mst5_rdata[(DWID - 1):0])
    ,.rid(mst5_rid[(IDWID - 1):0])
    ,.rlast(mst5_rlast)
    ,.rready(mst5_rready)
    ,.rresp(mst5_rresp[1:0])
    ,.rvalid(mst5_rvalid)
    ,.wdata(mst5_wdata[(DWID - 1):0])
    ,.wlast(mst5_wlast)
    ,.wready(mst5_wready)
    ,.wstrb(mst5_wstrb[(WSTRB - 1):0])
    ,.wvalid(mst5_wvalid)

    ,.a_araddr(split5_merge4_araddr[31:0])
    ,.a_arburst(split5_merge4_arburst[1:0])
    ,.a_arextras(split5_merge4_arextras[(EXTRAS - 1):0])
    ,.a_arid(split5_merge4_arid[(IDWID - 1):0])
    ,.a_arlen(split5_merge4_arlen[7:0])
    ,.a_arready(split5_merge4_arready)
    ,.a_arvalid(split5_merge4_arvalid)
    ,.a_awaddr(split5_merge4_awaddr[31:0])
    ,.a_awburst(split5_merge4_awburst[1:0])
    ,.a_awextras(split5_merge4_awextras[(EXTRAS - 1):0])
    ,.a_awid(split5_merge4_awid[(IDWID - 1):0])
    ,.a_awlen(split5_merge4_awlen[7:0])
    ,.a_awready(split5_merge4_awready)
    ,.a_awvalid(split5_merge4_awvalid)
    ,.a_bid(split5_merge4_bid[(IDWID - 1):0])
    ,.a_bready(split5_merge4_bready)
    ,.a_bresp(split5_merge4_bresp[1:0])
    ,.a_bvalid(split5_merge4_bvalid)
    ,.a_rdata(split5_merge4_rdata[(DWID - 1):0])
    ,.a_rid(split5_merge4_rid[(IDWID - 1):0])
    ,.a_rlast(split5_merge4_rlast)
    ,.a_rready(split5_merge4_rready)
    ,.a_rresp(split5_merge4_rresp[1:0])
    ,.a_rvalid(split5_merge4_rvalid)
    ,.a_wdata(split5_merge4_wdata[(DWID - 1):0])
    ,.a_wlast(split5_merge4_wlast)
    ,.a_wready(split5_merge4_wready)
    ,.a_wstrb(split5_merge4_wstrb[(WSTRB - 1):0])
    ,.a_wvalid(split5_merge4_wvalid)
    ,.b_araddr(split5_merge5_araddr[31:0])
    ,.b_arburst(split5_merge5_arburst[1:0])
    ,.b_arextras(split5_merge5_arextras[(EXTRAS - 1):0])
    ,.b_arid(split5_merge5_arid[(IDWID - 1):0])
    ,.b_arlen(split5_merge5_arlen[7:0])
    ,.b_arready(split5_merge5_arready)
    ,.b_arvalid(split5_merge5_arvalid)
    ,.b_awaddr(split5_merge5_awaddr[31:0])
    ,.b_awburst(split5_merge5_awburst[1:0])
    ,.b_awextras(split5_merge5_awextras[(EXTRAS - 1):0])
    ,.b_awid(split5_merge5_awid[(IDWID - 1):0])
    ,.b_awlen(split5_merge5_awlen[7:0])
    ,.b_awready(split5_merge5_awready)
    ,.b_awvalid(split5_merge5_awvalid)
    ,.b_bid(split5_merge5_bid[(IDWID - 1):0])
    ,.b_bready(split5_merge5_bready)
    ,.b_bresp(split5_merge5_bresp[1:0])
    ,.b_bvalid(split5_merge5_bvalid)
    ,.b_rdata(split5_merge5_rdata[(DWID - 1):0])
    ,.b_rid(split5_merge5_rid[(IDWID - 1):0])
    ,.b_rlast(split5_merge5_rlast)
    ,.b_rready(split5_merge5_rready)
    ,.b_rresp(split5_merge5_rresp[1:0])
    ,.b_rvalid(split5_merge5_rvalid)
    ,.b_wdata(split5_merge5_wdata[(DWID - 1):0])
    ,.b_wlast(split5_merge5_wlast)
    ,.b_wready(split5_merge5_wready)
    ,.b_wstrb(split5_merge5_wstrb[(WSTRB - 1):0])
    ,.b_wvalid(split5_merge5_wvalid)
    ,.c_araddr(split5_merge6_araddr[31:0])
    ,.c_arburst(split5_merge6_arburst[1:0])
    ,.c_arextras(split5_merge6_arextras[(EXTRAS - 1):0])
    ,.c_arid(split5_merge6_arid[(IDWID - 1):0])
    ,.c_arlen(split5_merge6_arlen[7:0])
    ,.c_arready(split5_merge6_arready)
    ,.c_arvalid(split5_merge6_arvalid)
    ,.c_awaddr(split5_merge6_awaddr[31:0])
    ,.c_awburst(split5_merge6_awburst[1:0])
    ,.c_awextras(split5_merge6_awextras[(EXTRAS - 1):0])
    ,.c_awid(split5_merge6_awid[(IDWID - 1):0])
    ,.c_awlen(split5_merge6_awlen[7:0])
    ,.c_awready(split5_merge6_awready)
    ,.c_awvalid(split5_merge6_awvalid)
    ,.c_bid(split5_merge6_bid[(IDWID - 1):0])
    ,.c_bready(split5_merge6_bready)
    ,.c_bresp(split5_merge6_bresp[1:0])
    ,.c_bvalid(split5_merge6_bvalid)
    ,.c_rdata(split5_merge6_rdata[(DWID - 1):0])
    ,.c_rid(split5_merge6_rid[(IDWID - 1):0])
    ,.c_rlast(split5_merge6_rlast)
    ,.c_rready(split5_merge6_rready)
    ,.c_rresp(split5_merge6_rresp[1:0])
    ,.c_rvalid(split5_merge6_rvalid)
    ,.c_wdata(split5_merge6_wdata[(DWID - 1):0])
    ,.c_wlast(split5_merge6_wlast)
    ,.c_wready(split5_merge6_wready)
    ,.c_wstrb(split5_merge6_wstrb[(WSTRB - 1):0])
    ,.c_wvalid(split5_merge6_wvalid)
    ,.d_araddr(split5_merge7_araddr[31:0])
    ,.d_arburst(split5_merge7_arburst[1:0])
    ,.d_arextras(split5_merge7_arextras[(EXTRAS - 1):0])
    ,.d_arid(split5_merge7_arid[(IDWID - 1):0])
    ,.d_arlen(split5_merge7_arlen[7:0])
    ,.d_arready(split5_merge7_arready)
    ,.d_arvalid(split5_merge7_arvalid)
    ,.d_awaddr(split5_merge7_awaddr[31:0])
    ,.d_awburst(split5_merge7_awburst[1:0])
    ,.d_awextras(split5_merge7_awextras[(EXTRAS - 1):0])
    ,.d_awid(split5_merge7_awid[(IDWID - 1):0])
    ,.d_awlen(split5_merge7_awlen[7:0])
    ,.d_awready(split5_merge7_awready)
    ,.d_awvalid(split5_merge7_awvalid)
    ,.d_bid(split5_merge7_bid[(IDWID - 1):0])
    ,.d_bready(split5_merge7_bready)
    ,.d_bresp(split5_merge7_bresp[1:0])
    ,.d_bvalid(split5_merge7_bvalid)
    ,.d_rdata(split5_merge7_rdata[(DWID - 1):0])
    ,.d_rid(split5_merge7_rid[(IDWID - 1):0])
    ,.d_rlast(split5_merge7_rlast)
    ,.d_rready(split5_merge7_rready)
    ,.d_rresp(split5_merge7_rresp[1:0])
    ,.d_rvalid(split5_merge7_rvalid)
    ,.d_wdata(split5_merge7_wdata[(DWID - 1):0])
    ,.d_wlast(split5_merge7_wlast)
    ,.d_wready(split5_merge7_wready)
    ,.d_wstrb(split5_merge7_wstrb[(WSTRB - 1):0])
    ,.d_wvalid(split5_merge7_wvalid)

);

axi_4_splitter split6 (
     .clk(clk) ,.rst_n(rst_n)

    ,.araddr(mst6_araddr[31:0])
    ,.arburst(mst6_arburst[1:0])
    ,.arextras(mst6_arextras[(EXTRAS - 1):0])
    ,.arid(mst6_arid[(IDWID - 1):0])
    ,.arlen(mst6_arlen[7:0])
    ,.arready(mst6_arready)
    ,.arvalid(mst6_arvalid)
    ,.awaddr(mst6_awaddr[31:0])
    ,.awburst(mst6_awburst[1:0])
    ,.awextras(mst6_awextras[(EXTRAS - 1):0])
    ,.awid(mst6_awid[3:0])
    ,.awlen(mst6_awlen[7:0])
    ,.awready(mst6_awready)
    ,.awvalid(mst6_awvalid)
    ,.bid(mst6_bid[(IDWID - 1):0])
    ,.bready(mst6_bready)
    ,.bresp(mst6_bresp[1:0])
    ,.bvalid(mst6_bvalid)
    ,.rdata(mst6_rdata[(DWID - 1):0])
    ,.rid(mst6_rid[(IDWID - 1):0])
    ,.rlast(mst6_rlast)
    ,.rready(mst6_rready)
    ,.rresp(mst6_rresp[1:0])
    ,.rvalid(mst6_rvalid)
    ,.wdata(mst6_wdata[(DWID - 1):0])
    ,.wlast(mst6_wlast)
    ,.wready(mst6_wready)
    ,.wstrb(mst6_wstrb[(WSTRB - 1):0])
    ,.wvalid(mst6_wvalid)

    ,.a_araddr(split6_merge4_araddr[31:0])
    ,.a_arburst(split6_merge4_arburst[1:0])
    ,.a_arextras(split6_merge4_arextras[(EXTRAS - 1):0])
    ,.a_arid(split6_merge4_arid[(IDWID - 1):0])
    ,.a_arlen(split6_merge4_arlen[7:0])
    ,.a_arready(split6_merge4_arready)
    ,.a_arvalid(split6_merge4_arvalid)
    ,.a_awaddr(split6_merge4_awaddr[31:0])
    ,.a_awburst(split6_merge4_awburst[1:0])
    ,.a_awextras(split6_merge4_awextras[(EXTRAS - 1):0])
    ,.a_awid(split6_merge4_awid[(IDWID - 1):0])
    ,.a_awlen(split6_merge4_awlen[7:0])
    ,.a_awready(split6_merge4_awready)
    ,.a_awvalid(split6_merge4_awvalid)
    ,.a_bid(split6_merge4_bid[(IDWID - 1):0])
    ,.a_bready(split6_merge4_bready)
    ,.a_bresp(split6_merge4_bresp[1:0])
    ,.a_bvalid(split6_merge4_bvalid)
    ,.a_rdata(split6_merge4_rdata[(DWID - 1):0])
    ,.a_rid(split6_merge4_rid[(IDWID - 1):0])
    ,.a_rlast(split6_merge4_rlast)
    ,.a_rready(split6_merge4_rready)
    ,.a_rresp(split6_merge4_rresp[1:0])
    ,.a_rvalid(split6_merge4_rvalid)
    ,.a_wdata(split6_merge4_wdata[(DWID - 1):0])
    ,.a_wlast(split6_merge4_wlast)
    ,.a_wready(split6_merge4_wready)
    ,.a_wstrb(split6_merge4_wstrb[(WSTRB - 1):0])
    ,.a_wvalid(split6_merge4_wvalid)
    ,.b_araddr(split6_merge5_araddr[31:0])
    ,.b_arburst(split6_merge5_arburst[1:0])
    ,.b_arextras(split6_merge5_arextras[(EXTRAS - 1):0])
    ,.b_arid(split6_merge5_arid[(IDWID - 1):0])
    ,.b_arlen(split6_merge5_arlen[7:0])
    ,.b_arready(split6_merge5_arready)
    ,.b_arvalid(split6_merge5_arvalid)
    ,.b_awaddr(split6_merge5_awaddr[31:0])
    ,.b_awburst(split6_merge5_awburst[1:0])
    ,.b_awextras(split6_merge5_awextras[(EXTRAS - 1):0])
    ,.b_awid(split6_merge5_awid[(IDWID - 1):0])
    ,.b_awlen(split6_merge5_awlen[7:0])
    ,.b_awready(split6_merge5_awready)
    ,.b_awvalid(split6_merge5_awvalid)
    ,.b_bid(split6_merge5_bid[(IDWID - 1):0])
    ,.b_bready(split6_merge5_bready)
    ,.b_bresp(split6_merge5_bresp[1:0])
    ,.b_bvalid(split6_merge5_bvalid)
    ,.b_rdata(split6_merge5_rdata[(DWID - 1):0])
    ,.b_rid(split6_merge5_rid[(IDWID - 1):0])
    ,.b_rlast(split6_merge5_rlast)
    ,.b_rready(split6_merge5_rready)
    ,.b_rresp(split6_merge5_rresp[1:0])
    ,.b_rvalid(split6_merge5_rvalid)
    ,.b_wdata(split6_merge5_wdata[(DWID - 1):0])
    ,.b_wlast(split6_merge5_wlast)
    ,.b_wready(split6_merge5_wready)
    ,.b_wstrb(split6_merge5_wstrb[(WSTRB - 1):0])
    ,.b_wvalid(split6_merge5_wvalid)
    ,.c_araddr(split6_merge6_araddr[31:0])
    ,.c_arburst(split6_merge6_arburst[1:0])
    ,.c_arextras(split6_merge6_arextras[(EXTRAS - 1):0])
    ,.c_arid(split6_merge6_arid[(IDWID - 1):0])
    ,.c_arlen(split6_merge6_arlen[7:0])
    ,.c_arready(split6_merge6_arready)
    ,.c_arvalid(split6_merge6_arvalid)
    ,.c_awaddr(split6_merge6_awaddr[31:0])
    ,.c_awburst(split6_merge6_awburst[1:0])
    ,.c_awextras(split6_merge6_awextras[(EXTRAS - 1):0])
    ,.c_awid(split6_merge6_awid[(IDWID - 1):0])
    ,.c_awlen(split6_merge6_awlen[7:0])
    ,.c_awready(split6_merge6_awready)
    ,.c_awvalid(split6_merge6_awvalid)
    ,.c_bid(split6_merge6_bid[(IDWID - 1):0])
    ,.c_bready(split6_merge6_bready)
    ,.c_bresp(split6_merge6_bresp[1:0])
    ,.c_bvalid(split6_merge6_bvalid)
    ,.c_rdata(split6_merge6_rdata[(DWID - 1):0])
    ,.c_rid(split6_merge6_rid[(IDWID - 1):0])
    ,.c_rlast(split6_merge6_rlast)
    ,.c_rready(split6_merge6_rready)
    ,.c_rresp(split6_merge6_rresp[1:0])
    ,.c_rvalid(split6_merge6_rvalid)
    ,.c_wdata(split6_merge6_wdata[(DWID - 1):0])
    ,.c_wlast(split6_merge6_wlast)
    ,.c_wready(split6_merge6_wready)
    ,.c_wstrb(split6_merge6_wstrb[(WSTRB - 1):0])
    ,.c_wvalid(split6_merge6_wvalid)
    ,.d_araddr(split6_merge7_araddr[31:0])
    ,.d_arburst(split6_merge7_arburst[1:0])
    ,.d_arextras(split6_merge7_arextras[(EXTRAS - 1):0])
    ,.d_arid(split6_merge7_arid[(IDWID - 1):0])
    ,.d_arlen(split6_merge7_arlen[7:0])
    ,.d_arready(split6_merge7_arready)
    ,.d_arvalid(split6_merge7_arvalid)
    ,.d_awaddr(split6_merge7_awaddr[31:0])
    ,.d_awburst(split6_merge7_awburst[1:0])
    ,.d_awextras(split6_merge7_awextras[(EXTRAS - 1):0])
    ,.d_awid(split6_merge7_awid[(IDWID - 1):0])
    ,.d_awlen(split6_merge7_awlen[7:0])
    ,.d_awready(split6_merge7_awready)
    ,.d_awvalid(split6_merge7_awvalid)
    ,.d_bid(split6_merge7_bid[(IDWID - 1):0])
    ,.d_bready(split6_merge7_bready)
    ,.d_bresp(split6_merge7_bresp[1:0])
    ,.d_bvalid(split6_merge7_bvalid)
    ,.d_rdata(split6_merge7_rdata[(DWID - 1):0])
    ,.d_rid(split6_merge7_rid[(IDWID - 1):0])
    ,.d_rlast(split6_merge7_rlast)
    ,.d_rready(split6_merge7_rready)
    ,.d_rresp(split6_merge7_rresp[1:0])
    ,.d_rvalid(split6_merge7_rvalid)
    ,.d_wdata(split6_merge7_wdata[(DWID - 1):0])
    ,.d_wlast(split6_merge7_wlast)
    ,.d_wready(split6_merge7_wready)
    ,.d_wstrb(split6_merge7_wstrb[(WSTRB - 1):0])
    ,.d_wvalid(split6_merge7_wvalid)

);

axi_4_splitter split7 (
     .clk(clk) ,.rst_n(rst_n)

    ,.araddr(mst7_araddr[31:0])
    ,.arburst(mst7_arburst[1:0])
    ,.arextras(mst7_arextras[(EXTRAS - 1):0])
    ,.arid(mst7_arid[(IDWID - 1):0])
    ,.arlen(mst7_arlen[7:0])
    ,.arready(mst7_arready)
    ,.arvalid(mst7_arvalid)
    ,.awaddr(mst7_awaddr[31:0])
    ,.awburst(mst7_awburst[1:0])
    ,.awextras(mst7_awextras[(EXTRAS - 1):0])
    ,.awid(mst7_awid[3:0])
    ,.awlen(mst7_awlen[7:0])
    ,.awready(mst7_awready)
    ,.awvalid(mst7_awvalid)
    ,.bid(mst7_bid[(IDWID - 1):0])
    ,.bready(mst7_bready)
    ,.bresp(mst7_bresp[1:0])
    ,.bvalid(mst7_bvalid)
    ,.rdata(mst7_rdata[(DWID - 1):0])
    ,.rid(mst7_rid[(IDWID - 1):0])
    ,.rlast(mst7_rlast)
    ,.rready(mst7_rready)
    ,.rresp(mst7_rresp[1:0])
    ,.rvalid(mst7_rvalid)
    ,.wdata(mst7_wdata[(DWID - 1):0])
    ,.wlast(mst7_wlast)
    ,.wready(mst7_wready)
    ,.wstrb(mst7_wstrb[(WSTRB - 1):0])
    ,.wvalid(mst7_wvalid)

    ,.a_araddr(split7_merge4_araddr[31:0])
    ,.a_arburst(split7_merge4_arburst[1:0])
    ,.a_arextras(split7_merge4_arextras[(EXTRAS - 1):0])
    ,.a_arid(split7_merge4_arid[(IDWID - 1):0])
    ,.a_arlen(split7_merge4_arlen[7:0])
    ,.a_arready(split7_merge4_arready)
    ,.a_arvalid(split7_merge4_arvalid)
    ,.a_awaddr(split7_merge4_awaddr[31:0])
    ,.a_awburst(split7_merge4_awburst[1:0])
    ,.a_awextras(split7_merge4_awextras[(EXTRAS - 1):0])
    ,.a_awid(split7_merge4_awid[(IDWID - 1):0])
    ,.a_awlen(split7_merge4_awlen[7:0])
    ,.a_awready(split7_merge4_awready)
    ,.a_awvalid(split7_merge4_awvalid)
    ,.a_bid(split7_merge4_bid[(IDWID - 1):0])
    ,.a_bready(split7_merge4_bready)
    ,.a_bresp(split7_merge4_bresp[1:0])
    ,.a_bvalid(split7_merge4_bvalid)
    ,.a_rdata(split7_merge4_rdata[(DWID - 1):0])
    ,.a_rid(split7_merge4_rid[(IDWID - 1):0])
    ,.a_rlast(split7_merge4_rlast)
    ,.a_rready(split7_merge4_rready)
    ,.a_rresp(split7_merge4_rresp[1:0])
    ,.a_rvalid(split7_merge4_rvalid)
    ,.a_wdata(split7_merge4_wdata[(DWID - 1):0])
    ,.a_wlast(split7_merge4_wlast)
    ,.a_wready(split7_merge4_wready)
    ,.a_wstrb(split7_merge4_wstrb[(WSTRB - 1):0])
    ,.a_wvalid(split7_merge4_wvalid)
    ,.b_araddr(split7_merge5_araddr[31:0])
    ,.b_arburst(split7_merge5_arburst[1:0])
    ,.b_arextras(split7_merge5_arextras[(EXTRAS - 1):0])
    ,.b_arid(split7_merge5_arid[(IDWID - 1):0])
    ,.b_arlen(split7_merge5_arlen[7:0])
    ,.b_arready(split7_merge5_arready)
    ,.b_arvalid(split7_merge5_arvalid)
    ,.b_awaddr(split7_merge5_awaddr[31:0])
    ,.b_awburst(split7_merge5_awburst[1:0])
    ,.b_awextras(split7_merge5_awextras[(EXTRAS - 1):0])
    ,.b_awid(split7_merge5_awid[(IDWID - 1):0])
    ,.b_awlen(split7_merge5_awlen[7:0])
    ,.b_awready(split7_merge5_awready)
    ,.b_awvalid(split7_merge5_awvalid)
    ,.b_bid(split7_merge5_bid[(IDWID - 1):0])
    ,.b_bready(split7_merge5_bready)
    ,.b_bresp(split7_merge5_bresp[1:0])
    ,.b_bvalid(split7_merge5_bvalid)
    ,.b_rdata(split7_merge5_rdata[(DWID - 1):0])
    ,.b_rid(split7_merge5_rid[(IDWID - 1):0])
    ,.b_rlast(split7_merge5_rlast)
    ,.b_rready(split7_merge5_rready)
    ,.b_rresp(split7_merge5_rresp[1:0])
    ,.b_rvalid(split7_merge5_rvalid)
    ,.b_wdata(split7_merge5_wdata[(DWID - 1):0])
    ,.b_wlast(split7_merge5_wlast)
    ,.b_wready(split7_merge5_wready)
    ,.b_wstrb(split7_merge5_wstrb[(WSTRB - 1):0])
    ,.b_wvalid(split7_merge5_wvalid)
    ,.c_araddr(split7_merge6_araddr[31:0])
    ,.c_arburst(split7_merge6_arburst[1:0])
    ,.c_arextras(split7_merge6_arextras[(EXTRAS - 1):0])
    ,.c_arid(split7_merge6_arid[(IDWID - 1):0])
    ,.c_arlen(split7_merge6_arlen[7:0])
    ,.c_arready(split7_merge6_arready)
    ,.c_arvalid(split7_merge6_arvalid)
    ,.c_awaddr(split7_merge6_awaddr[31:0])
    ,.c_awburst(split7_merge6_awburst[1:0])
    ,.c_awextras(split7_merge6_awextras[(EXTRAS - 1):0])
    ,.c_awid(split7_merge6_awid[(IDWID - 1):0])
    ,.c_awlen(split7_merge6_awlen[7:0])
    ,.c_awready(split7_merge6_awready)
    ,.c_awvalid(split7_merge6_awvalid)
    ,.c_bid(split7_merge6_bid[(IDWID - 1):0])
    ,.c_bready(split7_merge6_bready)
    ,.c_bresp(split7_merge6_bresp[1:0])
    ,.c_bvalid(split7_merge6_bvalid)
    ,.c_rdata(split7_merge6_rdata[(DWID - 1):0])
    ,.c_rid(split7_merge6_rid[(IDWID - 1):0])
    ,.c_rlast(split7_merge6_rlast)
    ,.c_rready(split7_merge6_rready)
    ,.c_rresp(split7_merge6_rresp[1:0])
    ,.c_rvalid(split7_merge6_rvalid)
    ,.c_wdata(split7_merge6_wdata[(DWID - 1):0])
    ,.c_wlast(split7_merge6_wlast)
    ,.c_wready(split7_merge6_wready)
    ,.c_wstrb(split7_merge6_wstrb[(WSTRB - 1):0])
    ,.c_wvalid(split7_merge6_wvalid)
    ,.d_araddr(split7_merge7_araddr[31:0])
    ,.d_arburst(split7_merge7_arburst[1:0])
    ,.d_arextras(split7_merge7_arextras[(EXTRAS - 1):0])
    ,.d_arid(split7_merge7_arid[(IDWID - 1):0])
    ,.d_arlen(split7_merge7_arlen[7:0])
    ,.d_arready(split7_merge7_arready)
    ,.d_arvalid(split7_merge7_arvalid)
    ,.d_awaddr(split7_merge7_awaddr[31:0])
    ,.d_awburst(split7_merge7_awburst[1:0])
    ,.d_awextras(split7_merge7_awextras[(EXTRAS - 1):0])
    ,.d_awid(split7_merge7_awid[(IDWID - 1):0])
    ,.d_awlen(split7_merge7_awlen[7:0])
    ,.d_awready(split7_merge7_awready)
    ,.d_awvalid(split7_merge7_awvalid)
    ,.d_bid(split7_merge7_bid[(IDWID - 1):0])
    ,.d_bready(split7_merge7_bready)
    ,.d_bresp(split7_merge7_bresp[1:0])
    ,.d_bvalid(split7_merge7_bvalid)
    ,.d_rdata(split7_merge7_rdata[(DWID - 1):0])
    ,.d_rid(split7_merge7_rid[(IDWID - 1):0])
    ,.d_rlast(split7_merge7_rlast)
    ,.d_rready(split7_merge7_rready)
    ,.d_rresp(split7_merge7_rresp[1:0])
    ,.d_rvalid(split7_merge7_rvalid)
    ,.d_wdata(split7_merge7_wdata[(DWID - 1):0])
    ,.d_wlast(split7_merge7_wlast)
    ,.d_wready(split7_merge7_wready)
    ,.d_wstrb(split7_merge7_wstrb[(WSTRB - 1):0])
    ,.d_wvalid(split7_merge7_wvalid)

);

wire [IDWID-1:0] split8_merge8_arid ;
wire [31:0] split8_merge8_araddr ;
wire [7:0] split8_merge8_arlen ;
wire [EXTRAS-1:0] split8_merge8_arextras ;
wire [1:0] split8_merge8_arburst ;
wire split8_merge8_arvalid ;
wire split8_merge8_arready ;
wire [IDWID-1:0] split8_merge8_rid ;
wire [DWID-1:0] split8_merge8_rdata ;
wire [1:0] split8_merge8_rresp ;
wire split8_merge8_rlast ;
wire split8_merge8_rvalid ;
wire split8_merge8_rready ;

wire [IDWID-1:0] split8_merge8_awid ;
wire [31:0] split8_merge8_awaddr ;
wire [7:0] split8_merge8_awlen ;
wire [EXTRAS-1:0] split8_merge8_awextras ;
wire [1:0] split8_merge8_awburst ;
wire split8_merge8_awvalid ;
wire split8_merge8_awready ;
wire [DWID-1:0] split8_merge8_wdata ;
wire [WSTRB-1:0] split8_merge8_wstrb ;
wire split8_merge8_wlast ;
wire split8_merge8_wvalid ;
wire split8_merge8_wready ;
wire [IDWID-1:0] split8_merge8_bid ;
wire [1:0] split8_merge8_bresp ;
wire split8_merge8_bvalid ;
wire split8_merge8_bready ;


wire [IDWID-1:0] split8_merge9_arid ;
wire [31:0] split8_merge9_araddr ;
wire [7:0] split8_merge9_arlen ;
wire [EXTRAS-1:0] split8_merge9_arextras ;
wire [1:0] split8_merge9_arburst ;
wire split8_merge9_arvalid ;
wire split8_merge9_arready ;
wire [IDWID-1:0] split8_merge9_rid ;
wire [DWID-1:0] split8_merge9_rdata ;
wire [1:0] split8_merge9_rresp ;
wire split8_merge9_rlast ;
wire split8_merge9_rvalid ;
wire split8_merge9_rready ;

wire [IDWID-1:0] split8_merge9_awid ;
wire [31:0] split8_merge9_awaddr ;
wire [7:0] split8_merge9_awlen ;
wire [EXTRAS-1:0] split8_merge9_awextras ;
wire [1:0] split8_merge9_awburst ;
wire split8_merge9_awvalid ;
wire split8_merge9_awready ;
wire [DWID-1:0] split8_merge9_wdata ;
wire [WSTRB-1:0] split8_merge9_wstrb ;
wire split8_merge9_wlast ;
wire split8_merge9_wvalid ;
wire split8_merge9_wready ;
wire [IDWID-1:0] split8_merge9_bid ;
wire [1:0] split8_merge9_bresp ;
wire split8_merge9_bvalid ;
wire split8_merge9_bready ;


wire [IDWID-1:0] split8_merge10_arid ;
wire [31:0] split8_merge10_araddr ;
wire [7:0] split8_merge10_arlen ;
wire [EXTRAS-1:0] split8_merge10_arextras ;
wire [1:0] split8_merge10_arburst ;
wire split8_merge10_arvalid ;
wire split8_merge10_arready ;
wire [IDWID-1:0] split8_merge10_rid ;
wire [DWID-1:0] split8_merge10_rdata ;
wire [1:0] split8_merge10_rresp ;
wire split8_merge10_rlast ;
wire split8_merge10_rvalid ;
wire split8_merge10_rready ;

wire [IDWID-1:0] split8_merge10_awid ;
wire [31:0] split8_merge10_awaddr ;
wire [7:0] split8_merge10_awlen ;
wire [EXTRAS-1:0] split8_merge10_awextras ;
wire [1:0] split8_merge10_awburst ;
wire split8_merge10_awvalid ;
wire split8_merge10_awready ;
wire [DWID-1:0] split8_merge10_wdata ;
wire [WSTRB-1:0] split8_merge10_wstrb ;
wire split8_merge10_wlast ;
wire split8_merge10_wvalid ;
wire split8_merge10_wready ;
wire [IDWID-1:0] split8_merge10_bid ;
wire [1:0] split8_merge10_bresp ;
wire split8_merge10_bvalid ;
wire split8_merge10_bready ;


wire [IDWID-1:0] split8_merge11_arid ;
wire [31:0] split8_merge11_araddr ;
wire [7:0] split8_merge11_arlen ;
wire [EXTRAS-1:0] split8_merge11_arextras ;
wire [1:0] split8_merge11_arburst ;
wire split8_merge11_arvalid ;
wire split8_merge11_arready ;
wire [IDWID-1:0] split8_merge11_rid ;
wire [DWID-1:0] split8_merge11_rdata ;
wire [1:0] split8_merge11_rresp ;
wire split8_merge11_rlast ;
wire split8_merge11_rvalid ;
wire split8_merge11_rready ;

wire [IDWID-1:0] split8_merge11_awid ;
wire [31:0] split8_merge11_awaddr ;
wire [7:0] split8_merge11_awlen ;
wire [EXTRAS-1:0] split8_merge11_awextras ;
wire [1:0] split8_merge11_awburst ;
wire split8_merge11_awvalid ;
wire split8_merge11_awready ;
wire [DWID-1:0] split8_merge11_wdata ;
wire [WSTRB-1:0] split8_merge11_wstrb ;
wire split8_merge11_wlast ;
wire split8_merge11_wvalid ;
wire split8_merge11_wready ;
wire [IDWID-1:0] split8_merge11_bid ;
wire [1:0] split8_merge11_bresp ;
wire split8_merge11_bvalid ;
wire split8_merge11_bready ;


axi_4_splitter split8 (
     .clk(clk) ,.rst_n(rst_n)

    ,.araddr(mst8_araddr[31:0])
    ,.arburst(mst8_arburst[1:0])
    ,.arextras(mst8_arextras[(EXTRAS - 1):0])
    ,.arid(mst8_arid[(IDWID - 1):0])
    ,.arlen(mst8_arlen[7:0])
    ,.arready(mst8_arready)
    ,.arvalid(mst8_arvalid)
    ,.awaddr(mst8_awaddr[31:0])
    ,.awburst(mst8_awburst[1:0])
    ,.awextras(mst8_awextras[(EXTRAS - 1):0])
    ,.awid(mst8_awid[3:0])
    ,.awlen(mst8_awlen[7:0])
    ,.awready(mst8_awready)
    ,.awvalid(mst8_awvalid)
    ,.bid(mst8_bid[(IDWID - 1):0])
    ,.bready(mst8_bready)
    ,.bresp(mst8_bresp[1:0])
    ,.bvalid(mst8_bvalid)
    ,.rdata(mst8_rdata[(DWID - 1):0])
    ,.rid(mst8_rid[(IDWID - 1):0])
    ,.rlast(mst8_rlast)
    ,.rready(mst8_rready)
    ,.rresp(mst8_rresp[1:0])
    ,.rvalid(mst8_rvalid)
    ,.wdata(mst8_wdata[(DWID - 1):0])
    ,.wlast(mst8_wlast)
    ,.wready(mst8_wready)
    ,.wstrb(mst8_wstrb[(WSTRB - 1):0])
    ,.wvalid(mst8_wvalid)

    ,.a_araddr(split8_merge8_araddr[31:0])
    ,.a_arburst(split8_merge8_arburst[1:0])
    ,.a_arextras(split8_merge8_arextras[(EXTRAS - 1):0])
    ,.a_arid(split8_merge8_arid[(IDWID - 1):0])
    ,.a_arlen(split8_merge8_arlen[7:0])
    ,.a_arready(split8_merge8_arready)
    ,.a_arvalid(split8_merge8_arvalid)
    ,.a_awaddr(split8_merge8_awaddr[31:0])
    ,.a_awburst(split8_merge8_awburst[1:0])
    ,.a_awextras(split8_merge8_awextras[(EXTRAS - 1):0])
    ,.a_awid(split8_merge8_awid[(IDWID - 1):0])
    ,.a_awlen(split8_merge8_awlen[7:0])
    ,.a_awready(split8_merge8_awready)
    ,.a_awvalid(split8_merge8_awvalid)
    ,.a_bid(split8_merge8_bid[(IDWID - 1):0])
    ,.a_bready(split8_merge8_bready)
    ,.a_bresp(split8_merge8_bresp[1:0])
    ,.a_bvalid(split8_merge8_bvalid)
    ,.a_rdata(split8_merge8_rdata[(DWID - 1):0])
    ,.a_rid(split8_merge8_rid[(IDWID - 1):0])
    ,.a_rlast(split8_merge8_rlast)
    ,.a_rready(split8_merge8_rready)
    ,.a_rresp(split8_merge8_rresp[1:0])
    ,.a_rvalid(split8_merge8_rvalid)
    ,.a_wdata(split8_merge8_wdata[(DWID - 1):0])
    ,.a_wlast(split8_merge8_wlast)
    ,.a_wready(split8_merge8_wready)
    ,.a_wstrb(split8_merge8_wstrb[(WSTRB - 1):0])
    ,.a_wvalid(split8_merge8_wvalid)
    ,.b_araddr(split8_merge9_araddr[31:0])
    ,.b_arburst(split8_merge9_arburst[1:0])
    ,.b_arextras(split8_merge9_arextras[(EXTRAS - 1):0])
    ,.b_arid(split8_merge9_arid[(IDWID - 1):0])
    ,.b_arlen(split8_merge9_arlen[7:0])
    ,.b_arready(split8_merge9_arready)
    ,.b_arvalid(split8_merge9_arvalid)
    ,.b_awaddr(split8_merge9_awaddr[31:0])
    ,.b_awburst(split8_merge9_awburst[1:0])
    ,.b_awextras(split8_merge9_awextras[(EXTRAS - 1):0])
    ,.b_awid(split8_merge9_awid[(IDWID - 1):0])
    ,.b_awlen(split8_merge9_awlen[7:0])
    ,.b_awready(split8_merge9_awready)
    ,.b_awvalid(split8_merge9_awvalid)
    ,.b_bid(split8_merge9_bid[(IDWID - 1):0])
    ,.b_bready(split8_merge9_bready)
    ,.b_bresp(split8_merge9_bresp[1:0])
    ,.b_bvalid(split8_merge9_bvalid)
    ,.b_rdata(split8_merge9_rdata[(DWID - 1):0])
    ,.b_rid(split8_merge9_rid[(IDWID - 1):0])
    ,.b_rlast(split8_merge9_rlast)
    ,.b_rready(split8_merge9_rready)
    ,.b_rresp(split8_merge9_rresp[1:0])
    ,.b_rvalid(split8_merge9_rvalid)
    ,.b_wdata(split8_merge9_wdata[(DWID - 1):0])
    ,.b_wlast(split8_merge9_wlast)
    ,.b_wready(split8_merge9_wready)
    ,.b_wstrb(split8_merge9_wstrb[(WSTRB - 1):0])
    ,.b_wvalid(split8_merge9_wvalid)
    ,.c_araddr(split8_merge10_araddr[31:0])
    ,.c_arburst(split8_merge10_arburst[1:0])
    ,.c_arextras(split8_merge10_arextras[(EXTRAS - 1):0])
    ,.c_arid(split8_merge10_arid[(IDWID - 1):0])
    ,.c_arlen(split8_merge10_arlen[7:0])
    ,.c_arready(split8_merge10_arready)
    ,.c_arvalid(split8_merge10_arvalid)
    ,.c_awaddr(split8_merge10_awaddr[31:0])
    ,.c_awburst(split8_merge10_awburst[1:0])
    ,.c_awextras(split8_merge10_awextras[(EXTRAS - 1):0])
    ,.c_awid(split8_merge10_awid[(IDWID - 1):0])
    ,.c_awlen(split8_merge10_awlen[7:0])
    ,.c_awready(split8_merge10_awready)
    ,.c_awvalid(split8_merge10_awvalid)
    ,.c_bid(split8_merge10_bid[(IDWID - 1):0])
    ,.c_bready(split8_merge10_bready)
    ,.c_bresp(split8_merge10_bresp[1:0])
    ,.c_bvalid(split8_merge10_bvalid)
    ,.c_rdata(split8_merge10_rdata[(DWID - 1):0])
    ,.c_rid(split8_merge10_rid[(IDWID - 1):0])
    ,.c_rlast(split8_merge10_rlast)
    ,.c_rready(split8_merge10_rready)
    ,.c_rresp(split8_merge10_rresp[1:0])
    ,.c_rvalid(split8_merge10_rvalid)
    ,.c_wdata(split8_merge10_wdata[(DWID - 1):0])
    ,.c_wlast(split8_merge10_wlast)
    ,.c_wready(split8_merge10_wready)
    ,.c_wstrb(split8_merge10_wstrb[(WSTRB - 1):0])
    ,.c_wvalid(split8_merge10_wvalid)
    ,.d_araddr(split8_merge11_araddr[31:0])
    ,.d_arburst(split8_merge11_arburst[1:0])
    ,.d_arextras(split8_merge11_arextras[(EXTRAS - 1):0])
    ,.d_arid(split8_merge11_arid[(IDWID - 1):0])
    ,.d_arlen(split8_merge11_arlen[7:0])
    ,.d_arready(split8_merge11_arready)
    ,.d_arvalid(split8_merge11_arvalid)
    ,.d_awaddr(split8_merge11_awaddr[31:0])
    ,.d_awburst(split8_merge11_awburst[1:0])
    ,.d_awextras(split8_merge11_awextras[(EXTRAS - 1):0])
    ,.d_awid(split8_merge11_awid[(IDWID - 1):0])
    ,.d_awlen(split8_merge11_awlen[7:0])
    ,.d_awready(split8_merge11_awready)
    ,.d_awvalid(split8_merge11_awvalid)
    ,.d_bid(split8_merge11_bid[(IDWID - 1):0])
    ,.d_bready(split8_merge11_bready)
    ,.d_bresp(split8_merge11_bresp[1:0])
    ,.d_bvalid(split8_merge11_bvalid)
    ,.d_rdata(split8_merge11_rdata[(DWID - 1):0])
    ,.d_rid(split8_merge11_rid[(IDWID - 1):0])
    ,.d_rlast(split8_merge11_rlast)
    ,.d_rready(split8_merge11_rready)
    ,.d_rresp(split8_merge11_rresp[1:0])
    ,.d_rvalid(split8_merge11_rvalid)
    ,.d_wdata(split8_merge11_wdata[(DWID - 1):0])
    ,.d_wlast(split8_merge11_wlast)
    ,.d_wready(split8_merge11_wready)
    ,.d_wstrb(split8_merge11_wstrb[(WSTRB - 1):0])
    ,.d_wvalid(split8_merge11_wvalid)

);

wire [IDWID-1:0] merge8_split108_arid ;
wire [31:0] merge8_split108_araddr ;
wire [7:0] merge8_split108_arlen ;
wire [EXTRAS-1:0] merge8_split108_arextras ;
wire [1:0] merge8_split108_arburst ;
wire merge8_split108_arvalid ;
wire merge8_split108_arready ;
wire [IDWID-1:0] merge8_split108_rid ;
wire [DWID-1:0] merge8_split108_rdata ;
wire [1:0] merge8_split108_rresp ;
wire merge8_split108_rlast ;
wire merge8_split108_rvalid ;
wire merge8_split108_rready ;

wire [IDWID-1:0] merge8_split108_awid ;
wire [31:0] merge8_split108_awaddr ;
wire [7:0] merge8_split108_awlen ;
wire [EXTRAS-1:0] merge8_split108_awextras ;
wire [1:0] merge8_split108_awburst ;
wire merge8_split108_awvalid ;
wire merge8_split108_awready ;
wire [DWID-1:0] merge8_split108_wdata ;
wire [WSTRB-1:0] merge8_split108_wstrb ;
wire merge8_split108_wlast ;
wire merge8_split108_wvalid ;
wire merge8_split108_wready ;
wire [IDWID-1:0] merge8_split108_bid ;
wire [1:0] merge8_split108_bresp ;
wire merge8_split108_bvalid ;
wire merge8_split108_bready ;


wire [IDWID-1:0] split9_merge8_arid ;
wire [31:0] split9_merge8_araddr ;
wire [7:0] split9_merge8_arlen ;
wire [EXTRAS-1:0] split9_merge8_arextras ;
wire [1:0] split9_merge8_arburst ;
wire split9_merge8_arvalid ;
wire split9_merge8_arready ;
wire [IDWID-1:0] split9_merge8_rid ;
wire [DWID-1:0] split9_merge8_rdata ;
wire [1:0] split9_merge8_rresp ;
wire split9_merge8_rlast ;
wire split9_merge8_rvalid ;
wire split9_merge8_rready ;

wire [IDWID-1:0] split9_merge8_awid ;
wire [31:0] split9_merge8_awaddr ;
wire [7:0] split9_merge8_awlen ;
wire [EXTRAS-1:0] split9_merge8_awextras ;
wire [1:0] split9_merge8_awburst ;
wire split9_merge8_awvalid ;
wire split9_merge8_awready ;
wire [DWID-1:0] split9_merge8_wdata ;
wire [WSTRB-1:0] split9_merge8_wstrb ;
wire split9_merge8_wlast ;
wire split9_merge8_wvalid ;
wire split9_merge8_wready ;
wire [IDWID-1:0] split9_merge8_bid ;
wire [1:0] split9_merge8_bresp ;
wire split9_merge8_bvalid ;
wire split9_merge8_bready ;


wire [IDWID-1:0] split10_merge8_arid ;
wire [31:0] split10_merge8_araddr ;
wire [7:0] split10_merge8_arlen ;
wire [EXTRAS-1:0] split10_merge8_arextras ;
wire [1:0] split10_merge8_arburst ;
wire split10_merge8_arvalid ;
wire split10_merge8_arready ;
wire [IDWID-1:0] split10_merge8_rid ;
wire [DWID-1:0] split10_merge8_rdata ;
wire [1:0] split10_merge8_rresp ;
wire split10_merge8_rlast ;
wire split10_merge8_rvalid ;
wire split10_merge8_rready ;

wire [IDWID-1:0] split10_merge8_awid ;
wire [31:0] split10_merge8_awaddr ;
wire [7:0] split10_merge8_awlen ;
wire [EXTRAS-1:0] split10_merge8_awextras ;
wire [1:0] split10_merge8_awburst ;
wire split10_merge8_awvalid ;
wire split10_merge8_awready ;
wire [DWID-1:0] split10_merge8_wdata ;
wire [WSTRB-1:0] split10_merge8_wstrb ;
wire split10_merge8_wlast ;
wire split10_merge8_wvalid ;
wire split10_merge8_wready ;
wire [IDWID-1:0] split10_merge8_bid ;
wire [1:0] split10_merge8_bresp ;
wire split10_merge8_bvalid ;
wire split10_merge8_bready ;


wire [IDWID-1:0] split11_merge8_arid ;
wire [31:0] split11_merge8_araddr ;
wire [7:0] split11_merge8_arlen ;
wire [EXTRAS-1:0] split11_merge8_arextras ;
wire [1:0] split11_merge8_arburst ;
wire split11_merge8_arvalid ;
wire split11_merge8_arready ;
wire [IDWID-1:0] split11_merge8_rid ;
wire [DWID-1:0] split11_merge8_rdata ;
wire [1:0] split11_merge8_rresp ;
wire split11_merge8_rlast ;
wire split11_merge8_rvalid ;
wire split11_merge8_rready ;

wire [IDWID-1:0] split11_merge8_awid ;
wire [31:0] split11_merge8_awaddr ;
wire [7:0] split11_merge8_awlen ;
wire [EXTRAS-1:0] split11_merge8_awextras ;
wire [1:0] split11_merge8_awburst ;
wire split11_merge8_awvalid ;
wire split11_merge8_awready ;
wire [DWID-1:0] split11_merge8_wdata ;
wire [WSTRB-1:0] split11_merge8_wstrb ;
wire split11_merge8_wlast ;
wire split11_merge8_wvalid ;
wire split11_merge8_wready ;
wire [IDWID-1:0] split11_merge8_bid ;
wire [1:0] split11_merge8_bresp ;
wire split11_merge8_bvalid ;
wire split11_merge8_bready ;


axi_4_merger merge8 (
     .clk(clk),.rst_n(rst_n)
    ,.araddr(merge8_split108_araddr[31:0])
    ,.arburst(merge8_split108_arburst[1:0])
    ,.arextras(merge8_split108_arextras[(EXTRAS - 1):0])
    ,.arid(merge8_split108_arid[(IDWID - 1):0])
    ,.arlen(merge8_split108_arlen[7:0])
    ,.arready(merge8_split108_arready)
    ,.arvalid(merge8_split108_arvalid)
    ,.awaddr(merge8_split108_awaddr[31:0])
    ,.awburst(merge8_split108_awburst[1:0])
    ,.awextras(merge8_split108_awextras[(EXTRAS - 1):0])
    ,.awid(merge8_split108_awid[3:0])
    ,.awlen(merge8_split108_awlen[7:0])
    ,.awready(merge8_split108_awready)
    ,.awvalid(merge8_split108_awvalid)
    ,.bid(merge8_split108_bid[(IDWID - 1):0])
    ,.bready(merge8_split108_bready)
    ,.bresp(merge8_split108_bresp[1:0])
    ,.bvalid(merge8_split108_bvalid)
    ,.rid(merge8_split108_rid[(IDWID - 1):0])
    ,.rlast(merge8_split108_rlast)
    ,.rready(merge8_split108_rready)
    ,.rresp(merge8_split108_rresp[1:0])
    ,.rvalid(merge8_split108_rvalid)
    ,.rdata(merge8_split108_rdata[(DWID - 1):0])
    ,.wdata(merge8_split108_wdata[(DWID - 1):0])
    ,.wlast(merge8_split108_wlast)
    ,.wready(merge8_split108_wready)
    ,.wstrb(merge8_split108_wstrb[(WSTRB - 1):0])
    ,.wvalid(merge8_split108_wvalid)


    ,.a_araddr(split8_merge8_araddr[31:0])
    ,.a_arburst(split8_merge8_arburst[1:0])
    ,.a_arextras(split8_merge8_arextras[(EXTRAS - 1):0])
    ,.a_arid(split8_merge8_arid[(IDWID - 1):0])
    ,.a_arlen(split8_merge8_arlen[7:0])
    ,.a_arready(split8_merge8_arready)
    ,.a_arvalid(split8_merge8_arvalid)
    ,.a_awaddr(split8_merge8_awaddr[31:0])
    ,.a_awburst(split8_merge8_awburst[1:0])
    ,.a_awextras(split8_merge8_awextras[(EXTRAS - 1):0])
    ,.a_awid(split8_merge8_awid[(IDWID - 1):0])
    ,.a_awlen(split8_merge8_awlen[7:0])
    ,.a_awready(split8_merge8_awready)
    ,.a_awvalid(split8_merge8_awvalid)
    ,.a_bid(split8_merge8_bid[(IDWID - 1):0])
    ,.a_bready(split8_merge8_bready)
    ,.a_bresp(split8_merge8_bresp[1:0])
    ,.a_bvalid(split8_merge8_bvalid)
    ,.a_rdata(split8_merge8_rdata[(DWID - 1):0])
    ,.a_rid(split8_merge8_rid[(IDWID - 1):0])
    ,.a_rlast(split8_merge8_rlast)
    ,.a_rready(split8_merge8_rready)
    ,.a_rresp(split8_merge8_rresp[1:0])
    ,.a_rvalid(split8_merge8_rvalid)
    ,.a_wdata(split8_merge8_wdata[(DWID - 1):0])
    ,.a_wlast(split8_merge8_wlast)
    ,.a_wready(split8_merge8_wready)
    ,.a_wstrb(split8_merge8_wstrb[(WSTRB - 1):0])
    ,.a_wvalid(split8_merge8_wvalid)

    ,.b_araddr(split9_merge8_araddr[31:0])
    ,.b_arburst(split9_merge8_arburst[1:0])
    ,.b_arextras(split9_merge8_arextras[(EXTRAS - 1):0])
    ,.b_arid(split9_merge8_arid[(IDWID - 1):0])
    ,.b_arlen(split9_merge8_arlen[7:0])
    ,.b_arready(split9_merge8_arready)
    ,.b_arvalid(split9_merge8_arvalid)
    ,.b_awaddr(split9_merge8_awaddr[31:0])
    ,.b_awburst(split9_merge8_awburst[1:0])
    ,.b_awextras(split9_merge8_awextras[(EXTRAS - 1):0])
    ,.b_awid(split9_merge8_awid[(IDWID - 1):0])
    ,.b_awlen(split9_merge8_awlen[7:0])
    ,.b_awready(split9_merge8_awready)
    ,.b_awvalid(split9_merge8_awvalid)
    ,.b_bid(split9_merge8_bid[(IDWID - 1):0])
    ,.b_bready(split9_merge8_bready)
    ,.b_bresp(split9_merge8_bresp[1:0])
    ,.b_bvalid(split9_merge8_bvalid)
    ,.b_rdata(split9_merge8_rdata[(DWID - 1):0])
    ,.b_rid(split9_merge8_rid[(IDWID - 1):0])
    ,.b_rlast(split9_merge8_rlast)
    ,.b_rready(split9_merge8_rready)
    ,.b_rresp(split9_merge8_rresp[1:0])
    ,.b_rvalid(split9_merge8_rvalid)
    ,.b_wdata(split9_merge8_wdata[(DWID - 1):0])
    ,.b_wlast(split9_merge8_wlast)
    ,.b_wready(split9_merge8_wready)
    ,.b_wstrb(split9_merge8_wstrb[(WSTRB - 1):0])
    ,.b_wvalid(split9_merge8_wvalid)

    ,.c_araddr(split10_merge8_araddr[31:0])
    ,.c_arburst(split10_merge8_arburst[1:0])
    ,.c_arextras(split10_merge8_arextras[(EXTRAS - 1):0])
    ,.c_arid(split10_merge8_arid[(IDWID - 1):0])
    ,.c_arlen(split10_merge8_arlen[7:0])
    ,.c_arready(split10_merge8_arready)
    ,.c_arvalid(split10_merge8_arvalid)
    ,.c_awaddr(split10_merge8_awaddr[31:0])
    ,.c_awburst(split10_merge8_awburst[1:0])
    ,.c_awextras(split10_merge8_awextras[(EXTRAS - 1):0])
    ,.c_awid(split10_merge8_awid[(IDWID - 1):0])
    ,.c_awlen(split10_merge8_awlen[7:0])
    ,.c_awready(split10_merge8_awready)
    ,.c_awvalid(split10_merge8_awvalid)
    ,.c_bid(split10_merge8_bid[(IDWID - 1):0])
    ,.c_bready(split10_merge8_bready)
    ,.c_bresp(split10_merge8_bresp[1:0])
    ,.c_bvalid(split10_merge8_bvalid)
    ,.c_rdata(split10_merge8_rdata[(DWID - 1):0])
    ,.c_rid(split10_merge8_rid[(IDWID - 1):0])
    ,.c_rlast(split10_merge8_rlast)
    ,.c_rready(split10_merge8_rready)
    ,.c_rresp(split10_merge8_rresp[1:0])
    ,.c_rvalid(split10_merge8_rvalid)
    ,.c_wdata(split10_merge8_wdata[(DWID - 1):0])
    ,.c_wlast(split10_merge8_wlast)
    ,.c_wready(split10_merge8_wready)
    ,.c_wstrb(split10_merge8_wstrb[(WSTRB - 1):0])
    ,.c_wvalid(split10_merge8_wvalid)

    ,.d_araddr(split11_merge8_araddr[31:0])
    ,.d_arburst(split11_merge8_arburst[1:0])
    ,.d_arextras(split11_merge8_arextras[(EXTRAS - 1):0])
    ,.d_arid(split11_merge8_arid[(IDWID - 1):0])
    ,.d_arlen(split11_merge8_arlen[7:0])
    ,.d_arready(split11_merge8_arready)
    ,.d_arvalid(split11_merge8_arvalid)
    ,.d_awaddr(split11_merge8_awaddr[31:0])
    ,.d_awburst(split11_merge8_awburst[1:0])
    ,.d_awextras(split11_merge8_awextras[(EXTRAS - 1):0])
    ,.d_awid(split11_merge8_awid[(IDWID - 1):0])
    ,.d_awlen(split11_merge8_awlen[7:0])
    ,.d_awready(split11_merge8_awready)
    ,.d_awvalid(split11_merge8_awvalid)
    ,.d_bid(split11_merge8_bid[(IDWID - 1):0])
    ,.d_bready(split11_merge8_bready)
    ,.d_bresp(split11_merge8_bresp[1:0])
    ,.d_bvalid(split11_merge8_bvalid)
    ,.d_rdata(split11_merge8_rdata[(DWID - 1):0])
    ,.d_rid(split11_merge8_rid[(IDWID - 1):0])
    ,.d_rlast(split11_merge8_rlast)
    ,.d_rready(split11_merge8_rready)
    ,.d_rresp(split11_merge8_rresp[1:0])
    ,.d_rvalid(split11_merge8_rvalid)
    ,.d_wdata(split11_merge8_wdata[(DWID - 1):0])
    ,.d_wlast(split11_merge8_wlast)
    ,.d_wready(split11_merge8_wready)
    ,.d_wstrb(split11_merge8_wstrb[(WSTRB - 1):0])
    ,.d_wvalid(split11_merge8_wvalid)
);


wire [IDWID-1:0] merge9_split109_arid ;
wire [31:0] merge9_split109_araddr ;
wire [7:0] merge9_split109_arlen ;
wire [EXTRAS-1:0] merge9_split109_arextras ;
wire [1:0] merge9_split109_arburst ;
wire merge9_split109_arvalid ;
wire merge9_split109_arready ;
wire [IDWID-1:0] merge9_split109_rid ;
wire [DWID-1:0] merge9_split109_rdata ;
wire [1:0] merge9_split109_rresp ;
wire merge9_split109_rlast ;
wire merge9_split109_rvalid ;
wire merge9_split109_rready ;

wire [IDWID-1:0] merge9_split109_awid ;
wire [31:0] merge9_split109_awaddr ;
wire [7:0] merge9_split109_awlen ;
wire [EXTRAS-1:0] merge9_split109_awextras ;
wire [1:0] merge9_split109_awburst ;
wire merge9_split109_awvalid ;
wire merge9_split109_awready ;
wire [DWID-1:0] merge9_split109_wdata ;
wire [WSTRB-1:0] merge9_split109_wstrb ;
wire merge9_split109_wlast ;
wire merge9_split109_wvalid ;
wire merge9_split109_wready ;
wire [IDWID-1:0] merge9_split109_bid ;
wire [1:0] merge9_split109_bresp ;
wire merge9_split109_bvalid ;
wire merge9_split109_bready ;


wire [IDWID-1:0] split9_merge9_arid ;
wire [31:0] split9_merge9_araddr ;
wire [7:0] split9_merge9_arlen ;
wire [EXTRAS-1:0] split9_merge9_arextras ;
wire [1:0] split9_merge9_arburst ;
wire split9_merge9_arvalid ;
wire split9_merge9_arready ;
wire [IDWID-1:0] split9_merge9_rid ;
wire [DWID-1:0] split9_merge9_rdata ;
wire [1:0] split9_merge9_rresp ;
wire split9_merge9_rlast ;
wire split9_merge9_rvalid ;
wire split9_merge9_rready ;

wire [IDWID-1:0] split9_merge9_awid ;
wire [31:0] split9_merge9_awaddr ;
wire [7:0] split9_merge9_awlen ;
wire [EXTRAS-1:0] split9_merge9_awextras ;
wire [1:0] split9_merge9_awburst ;
wire split9_merge9_awvalid ;
wire split9_merge9_awready ;
wire [DWID-1:0] split9_merge9_wdata ;
wire [WSTRB-1:0] split9_merge9_wstrb ;
wire split9_merge9_wlast ;
wire split9_merge9_wvalid ;
wire split9_merge9_wready ;
wire [IDWID-1:0] split9_merge9_bid ;
wire [1:0] split9_merge9_bresp ;
wire split9_merge9_bvalid ;
wire split9_merge9_bready ;


wire [IDWID-1:0] split10_merge9_arid ;
wire [31:0] split10_merge9_araddr ;
wire [7:0] split10_merge9_arlen ;
wire [EXTRAS-1:0] split10_merge9_arextras ;
wire [1:0] split10_merge9_arburst ;
wire split10_merge9_arvalid ;
wire split10_merge9_arready ;
wire [IDWID-1:0] split10_merge9_rid ;
wire [DWID-1:0] split10_merge9_rdata ;
wire [1:0] split10_merge9_rresp ;
wire split10_merge9_rlast ;
wire split10_merge9_rvalid ;
wire split10_merge9_rready ;

wire [IDWID-1:0] split10_merge9_awid ;
wire [31:0] split10_merge9_awaddr ;
wire [7:0] split10_merge9_awlen ;
wire [EXTRAS-1:0] split10_merge9_awextras ;
wire [1:0] split10_merge9_awburst ;
wire split10_merge9_awvalid ;
wire split10_merge9_awready ;
wire [DWID-1:0] split10_merge9_wdata ;
wire [WSTRB-1:0] split10_merge9_wstrb ;
wire split10_merge9_wlast ;
wire split10_merge9_wvalid ;
wire split10_merge9_wready ;
wire [IDWID-1:0] split10_merge9_bid ;
wire [1:0] split10_merge9_bresp ;
wire split10_merge9_bvalid ;
wire split10_merge9_bready ;


wire [IDWID-1:0] split11_merge9_arid ;
wire [31:0] split11_merge9_araddr ;
wire [7:0] split11_merge9_arlen ;
wire [EXTRAS-1:0] split11_merge9_arextras ;
wire [1:0] split11_merge9_arburst ;
wire split11_merge9_arvalid ;
wire split11_merge9_arready ;
wire [IDWID-1:0] split11_merge9_rid ;
wire [DWID-1:0] split11_merge9_rdata ;
wire [1:0] split11_merge9_rresp ;
wire split11_merge9_rlast ;
wire split11_merge9_rvalid ;
wire split11_merge9_rready ;

wire [IDWID-1:0] split11_merge9_awid ;
wire [31:0] split11_merge9_awaddr ;
wire [7:0] split11_merge9_awlen ;
wire [EXTRAS-1:0] split11_merge9_awextras ;
wire [1:0] split11_merge9_awburst ;
wire split11_merge9_awvalid ;
wire split11_merge9_awready ;
wire [DWID-1:0] split11_merge9_wdata ;
wire [WSTRB-1:0] split11_merge9_wstrb ;
wire split11_merge9_wlast ;
wire split11_merge9_wvalid ;
wire split11_merge9_wready ;
wire [IDWID-1:0] split11_merge9_bid ;
wire [1:0] split11_merge9_bresp ;
wire split11_merge9_bvalid ;
wire split11_merge9_bready ;


axi_4_merger merge9 (
     .clk(clk),.rst_n(rst_n)
    ,.araddr(merge9_split109_araddr[31:0])
    ,.arburst(merge9_split109_arburst[1:0])
    ,.arextras(merge9_split109_arextras[(EXTRAS - 1):0])
    ,.arid(merge9_split109_arid[(IDWID - 1):0])
    ,.arlen(merge9_split109_arlen[7:0])
    ,.arready(merge9_split109_arready)
    ,.arvalid(merge9_split109_arvalid)
    ,.awaddr(merge9_split109_awaddr[31:0])
    ,.awburst(merge9_split109_awburst[1:0])
    ,.awextras(merge9_split109_awextras[(EXTRAS - 1):0])
    ,.awid(merge9_split109_awid[3:0])
    ,.awlen(merge9_split109_awlen[7:0])
    ,.awready(merge9_split109_awready)
    ,.awvalid(merge9_split109_awvalid)
    ,.bid(merge9_split109_bid[(IDWID - 1):0])
    ,.bready(merge9_split109_bready)
    ,.bresp(merge9_split109_bresp[1:0])
    ,.bvalid(merge9_split109_bvalid)
    ,.rid(merge9_split109_rid[(IDWID - 1):0])
    ,.rlast(merge9_split109_rlast)
    ,.rready(merge9_split109_rready)
    ,.rresp(merge9_split109_rresp[1:0])
    ,.rvalid(merge9_split109_rvalid)
    ,.rdata(merge9_split109_rdata[(DWID - 1):0])
    ,.wdata(merge9_split109_wdata[(DWID - 1):0])
    ,.wlast(merge9_split109_wlast)
    ,.wready(merge9_split109_wready)
    ,.wstrb(merge9_split109_wstrb[(WSTRB - 1):0])
    ,.wvalid(merge9_split109_wvalid)


    ,.a_araddr(split8_merge9_araddr[31:0])
    ,.a_arburst(split8_merge9_arburst[1:0])
    ,.a_arextras(split8_merge9_arextras[(EXTRAS - 1):0])
    ,.a_arid(split8_merge9_arid[(IDWID - 1):0])
    ,.a_arlen(split8_merge9_arlen[7:0])
    ,.a_arready(split8_merge9_arready)
    ,.a_arvalid(split8_merge9_arvalid)
    ,.a_awaddr(split8_merge9_awaddr[31:0])
    ,.a_awburst(split8_merge9_awburst[1:0])
    ,.a_awextras(split8_merge9_awextras[(EXTRAS - 1):0])
    ,.a_awid(split8_merge9_awid[(IDWID - 1):0])
    ,.a_awlen(split8_merge9_awlen[7:0])
    ,.a_awready(split8_merge9_awready)
    ,.a_awvalid(split8_merge9_awvalid)
    ,.a_bid(split8_merge9_bid[(IDWID - 1):0])
    ,.a_bready(split8_merge9_bready)
    ,.a_bresp(split8_merge9_bresp[1:0])
    ,.a_bvalid(split8_merge9_bvalid)
    ,.a_rdata(split8_merge9_rdata[(DWID - 1):0])
    ,.a_rid(split8_merge9_rid[(IDWID - 1):0])
    ,.a_rlast(split8_merge9_rlast)
    ,.a_rready(split8_merge9_rready)
    ,.a_rresp(split8_merge9_rresp[1:0])
    ,.a_rvalid(split8_merge9_rvalid)
    ,.a_wdata(split8_merge9_wdata[(DWID - 1):0])
    ,.a_wlast(split8_merge9_wlast)
    ,.a_wready(split8_merge9_wready)
    ,.a_wstrb(split8_merge9_wstrb[(WSTRB - 1):0])
    ,.a_wvalid(split8_merge9_wvalid)

    ,.b_araddr(split9_merge9_araddr[31:0])
    ,.b_arburst(split9_merge9_arburst[1:0])
    ,.b_arextras(split9_merge9_arextras[(EXTRAS - 1):0])
    ,.b_arid(split9_merge9_arid[(IDWID - 1):0])
    ,.b_arlen(split9_merge9_arlen[7:0])
    ,.b_arready(split9_merge9_arready)
    ,.b_arvalid(split9_merge9_arvalid)
    ,.b_awaddr(split9_merge9_awaddr[31:0])
    ,.b_awburst(split9_merge9_awburst[1:0])
    ,.b_awextras(split9_merge9_awextras[(EXTRAS - 1):0])
    ,.b_awid(split9_merge9_awid[(IDWID - 1):0])
    ,.b_awlen(split9_merge9_awlen[7:0])
    ,.b_awready(split9_merge9_awready)
    ,.b_awvalid(split9_merge9_awvalid)
    ,.b_bid(split9_merge9_bid[(IDWID - 1):0])
    ,.b_bready(split9_merge9_bready)
    ,.b_bresp(split9_merge9_bresp[1:0])
    ,.b_bvalid(split9_merge9_bvalid)
    ,.b_rdata(split9_merge9_rdata[(DWID - 1):0])
    ,.b_rid(split9_merge9_rid[(IDWID - 1):0])
    ,.b_rlast(split9_merge9_rlast)
    ,.b_rready(split9_merge9_rready)
    ,.b_rresp(split9_merge9_rresp[1:0])
    ,.b_rvalid(split9_merge9_rvalid)
    ,.b_wdata(split9_merge9_wdata[(DWID - 1):0])
    ,.b_wlast(split9_merge9_wlast)
    ,.b_wready(split9_merge9_wready)
    ,.b_wstrb(split9_merge9_wstrb[(WSTRB - 1):0])
    ,.b_wvalid(split9_merge9_wvalid)

    ,.c_araddr(split10_merge9_araddr[31:0])
    ,.c_arburst(split10_merge9_arburst[1:0])
    ,.c_arextras(split10_merge9_arextras[(EXTRAS - 1):0])
    ,.c_arid(split10_merge9_arid[(IDWID - 1):0])
    ,.c_arlen(split10_merge9_arlen[7:0])
    ,.c_arready(split10_merge9_arready)
    ,.c_arvalid(split10_merge9_arvalid)
    ,.c_awaddr(split10_merge9_awaddr[31:0])
    ,.c_awburst(split10_merge9_awburst[1:0])
    ,.c_awextras(split10_merge9_awextras[(EXTRAS - 1):0])
    ,.c_awid(split10_merge9_awid[(IDWID - 1):0])
    ,.c_awlen(split10_merge9_awlen[7:0])
    ,.c_awready(split10_merge9_awready)
    ,.c_awvalid(split10_merge9_awvalid)
    ,.c_bid(split10_merge9_bid[(IDWID - 1):0])
    ,.c_bready(split10_merge9_bready)
    ,.c_bresp(split10_merge9_bresp[1:0])
    ,.c_bvalid(split10_merge9_bvalid)
    ,.c_rdata(split10_merge9_rdata[(DWID - 1):0])
    ,.c_rid(split10_merge9_rid[(IDWID - 1):0])
    ,.c_rlast(split10_merge9_rlast)
    ,.c_rready(split10_merge9_rready)
    ,.c_rresp(split10_merge9_rresp[1:0])
    ,.c_rvalid(split10_merge9_rvalid)
    ,.c_wdata(split10_merge9_wdata[(DWID - 1):0])
    ,.c_wlast(split10_merge9_wlast)
    ,.c_wready(split10_merge9_wready)
    ,.c_wstrb(split10_merge9_wstrb[(WSTRB - 1):0])
    ,.c_wvalid(split10_merge9_wvalid)

    ,.d_araddr(split11_merge9_araddr[31:0])
    ,.d_arburst(split11_merge9_arburst[1:0])
    ,.d_arextras(split11_merge9_arextras[(EXTRAS - 1):0])
    ,.d_arid(split11_merge9_arid[(IDWID - 1):0])
    ,.d_arlen(split11_merge9_arlen[7:0])
    ,.d_arready(split11_merge9_arready)
    ,.d_arvalid(split11_merge9_arvalid)
    ,.d_awaddr(split11_merge9_awaddr[31:0])
    ,.d_awburst(split11_merge9_awburst[1:0])
    ,.d_awextras(split11_merge9_awextras[(EXTRAS - 1):0])
    ,.d_awid(split11_merge9_awid[(IDWID - 1):0])
    ,.d_awlen(split11_merge9_awlen[7:0])
    ,.d_awready(split11_merge9_awready)
    ,.d_awvalid(split11_merge9_awvalid)
    ,.d_bid(split11_merge9_bid[(IDWID - 1):0])
    ,.d_bready(split11_merge9_bready)
    ,.d_bresp(split11_merge9_bresp[1:0])
    ,.d_bvalid(split11_merge9_bvalid)
    ,.d_rdata(split11_merge9_rdata[(DWID - 1):0])
    ,.d_rid(split11_merge9_rid[(IDWID - 1):0])
    ,.d_rlast(split11_merge9_rlast)
    ,.d_rready(split11_merge9_rready)
    ,.d_rresp(split11_merge9_rresp[1:0])
    ,.d_rvalid(split11_merge9_rvalid)
    ,.d_wdata(split11_merge9_wdata[(DWID - 1):0])
    ,.d_wlast(split11_merge9_wlast)
    ,.d_wready(split11_merge9_wready)
    ,.d_wstrb(split11_merge9_wstrb[(WSTRB - 1):0])
    ,.d_wvalid(split11_merge9_wvalid)
);


wire [IDWID-1:0] merge10_split110_arid ;
wire [31:0] merge10_split110_araddr ;
wire [7:0] merge10_split110_arlen ;
wire [EXTRAS-1:0] merge10_split110_arextras ;
wire [1:0] merge10_split110_arburst ;
wire merge10_split110_arvalid ;
wire merge10_split110_arready ;
wire [IDWID-1:0] merge10_split110_rid ;
wire [DWID-1:0] merge10_split110_rdata ;
wire [1:0] merge10_split110_rresp ;
wire merge10_split110_rlast ;
wire merge10_split110_rvalid ;
wire merge10_split110_rready ;

wire [IDWID-1:0] merge10_split110_awid ;
wire [31:0] merge10_split110_awaddr ;
wire [7:0] merge10_split110_awlen ;
wire [EXTRAS-1:0] merge10_split110_awextras ;
wire [1:0] merge10_split110_awburst ;
wire merge10_split110_awvalid ;
wire merge10_split110_awready ;
wire [DWID-1:0] merge10_split110_wdata ;
wire [WSTRB-1:0] merge10_split110_wstrb ;
wire merge10_split110_wlast ;
wire merge10_split110_wvalid ;
wire merge10_split110_wready ;
wire [IDWID-1:0] merge10_split110_bid ;
wire [1:0] merge10_split110_bresp ;
wire merge10_split110_bvalid ;
wire merge10_split110_bready ;


wire [IDWID-1:0] split9_merge10_arid ;
wire [31:0] split9_merge10_araddr ;
wire [7:0] split9_merge10_arlen ;
wire [EXTRAS-1:0] split9_merge10_arextras ;
wire [1:0] split9_merge10_arburst ;
wire split9_merge10_arvalid ;
wire split9_merge10_arready ;
wire [IDWID-1:0] split9_merge10_rid ;
wire [DWID-1:0] split9_merge10_rdata ;
wire [1:0] split9_merge10_rresp ;
wire split9_merge10_rlast ;
wire split9_merge10_rvalid ;
wire split9_merge10_rready ;

wire [IDWID-1:0] split9_merge10_awid ;
wire [31:0] split9_merge10_awaddr ;
wire [7:0] split9_merge10_awlen ;
wire [EXTRAS-1:0] split9_merge10_awextras ;
wire [1:0] split9_merge10_awburst ;
wire split9_merge10_awvalid ;
wire split9_merge10_awready ;
wire [DWID-1:0] split9_merge10_wdata ;
wire [WSTRB-1:0] split9_merge10_wstrb ;
wire split9_merge10_wlast ;
wire split9_merge10_wvalid ;
wire split9_merge10_wready ;
wire [IDWID-1:0] split9_merge10_bid ;
wire [1:0] split9_merge10_bresp ;
wire split9_merge10_bvalid ;
wire split9_merge10_bready ;


wire [IDWID-1:0] split10_merge10_arid ;
wire [31:0] split10_merge10_araddr ;
wire [7:0] split10_merge10_arlen ;
wire [EXTRAS-1:0] split10_merge10_arextras ;
wire [1:0] split10_merge10_arburst ;
wire split10_merge10_arvalid ;
wire split10_merge10_arready ;
wire [IDWID-1:0] split10_merge10_rid ;
wire [DWID-1:0] split10_merge10_rdata ;
wire [1:0] split10_merge10_rresp ;
wire split10_merge10_rlast ;
wire split10_merge10_rvalid ;
wire split10_merge10_rready ;

wire [IDWID-1:0] split10_merge10_awid ;
wire [31:0] split10_merge10_awaddr ;
wire [7:0] split10_merge10_awlen ;
wire [EXTRAS-1:0] split10_merge10_awextras ;
wire [1:0] split10_merge10_awburst ;
wire split10_merge10_awvalid ;
wire split10_merge10_awready ;
wire [DWID-1:0] split10_merge10_wdata ;
wire [WSTRB-1:0] split10_merge10_wstrb ;
wire split10_merge10_wlast ;
wire split10_merge10_wvalid ;
wire split10_merge10_wready ;
wire [IDWID-1:0] split10_merge10_bid ;
wire [1:0] split10_merge10_bresp ;
wire split10_merge10_bvalid ;
wire split10_merge10_bready ;


wire [IDWID-1:0] split11_merge10_arid ;
wire [31:0] split11_merge10_araddr ;
wire [7:0] split11_merge10_arlen ;
wire [EXTRAS-1:0] split11_merge10_arextras ;
wire [1:0] split11_merge10_arburst ;
wire split11_merge10_arvalid ;
wire split11_merge10_arready ;
wire [IDWID-1:0] split11_merge10_rid ;
wire [DWID-1:0] split11_merge10_rdata ;
wire [1:0] split11_merge10_rresp ;
wire split11_merge10_rlast ;
wire split11_merge10_rvalid ;
wire split11_merge10_rready ;

wire [IDWID-1:0] split11_merge10_awid ;
wire [31:0] split11_merge10_awaddr ;
wire [7:0] split11_merge10_awlen ;
wire [EXTRAS-1:0] split11_merge10_awextras ;
wire [1:0] split11_merge10_awburst ;
wire split11_merge10_awvalid ;
wire split11_merge10_awready ;
wire [DWID-1:0] split11_merge10_wdata ;
wire [WSTRB-1:0] split11_merge10_wstrb ;
wire split11_merge10_wlast ;
wire split11_merge10_wvalid ;
wire split11_merge10_wready ;
wire [IDWID-1:0] split11_merge10_bid ;
wire [1:0] split11_merge10_bresp ;
wire split11_merge10_bvalid ;
wire split11_merge10_bready ;


axi_4_merger merge10 (
     .clk(clk),.rst_n(rst_n)
    ,.araddr(merge10_split110_araddr[31:0])
    ,.arburst(merge10_split110_arburst[1:0])
    ,.arextras(merge10_split110_arextras[(EXTRAS - 1):0])
    ,.arid(merge10_split110_arid[(IDWID - 1):0])
    ,.arlen(merge10_split110_arlen[7:0])
    ,.arready(merge10_split110_arready)
    ,.arvalid(merge10_split110_arvalid)
    ,.awaddr(merge10_split110_awaddr[31:0])
    ,.awburst(merge10_split110_awburst[1:0])
    ,.awextras(merge10_split110_awextras[(EXTRAS - 1):0])
    ,.awid(merge10_split110_awid[3:0])
    ,.awlen(merge10_split110_awlen[7:0])
    ,.awready(merge10_split110_awready)
    ,.awvalid(merge10_split110_awvalid)
    ,.bid(merge10_split110_bid[(IDWID - 1):0])
    ,.bready(merge10_split110_bready)
    ,.bresp(merge10_split110_bresp[1:0])
    ,.bvalid(merge10_split110_bvalid)
    ,.rid(merge10_split110_rid[(IDWID - 1):0])
    ,.rlast(merge10_split110_rlast)
    ,.rready(merge10_split110_rready)
    ,.rresp(merge10_split110_rresp[1:0])
    ,.rvalid(merge10_split110_rvalid)
    ,.rdata(merge10_split110_rdata[(DWID - 1):0])
    ,.wdata(merge10_split110_wdata[(DWID - 1):0])
    ,.wlast(merge10_split110_wlast)
    ,.wready(merge10_split110_wready)
    ,.wstrb(merge10_split110_wstrb[(WSTRB - 1):0])
    ,.wvalid(merge10_split110_wvalid)


    ,.a_araddr(split8_merge10_araddr[31:0])
    ,.a_arburst(split8_merge10_arburst[1:0])
    ,.a_arextras(split8_merge10_arextras[(EXTRAS - 1):0])
    ,.a_arid(split8_merge10_arid[(IDWID - 1):0])
    ,.a_arlen(split8_merge10_arlen[7:0])
    ,.a_arready(split8_merge10_arready)
    ,.a_arvalid(split8_merge10_arvalid)
    ,.a_awaddr(split8_merge10_awaddr[31:0])
    ,.a_awburst(split8_merge10_awburst[1:0])
    ,.a_awextras(split8_merge10_awextras[(EXTRAS - 1):0])
    ,.a_awid(split8_merge10_awid[(IDWID - 1):0])
    ,.a_awlen(split8_merge10_awlen[7:0])
    ,.a_awready(split8_merge10_awready)
    ,.a_awvalid(split8_merge10_awvalid)
    ,.a_bid(split8_merge10_bid[(IDWID - 1):0])
    ,.a_bready(split8_merge10_bready)
    ,.a_bresp(split8_merge10_bresp[1:0])
    ,.a_bvalid(split8_merge10_bvalid)
    ,.a_rdata(split8_merge10_rdata[(DWID - 1):0])
    ,.a_rid(split8_merge10_rid[(IDWID - 1):0])
    ,.a_rlast(split8_merge10_rlast)
    ,.a_rready(split8_merge10_rready)
    ,.a_rresp(split8_merge10_rresp[1:0])
    ,.a_rvalid(split8_merge10_rvalid)
    ,.a_wdata(split8_merge10_wdata[(DWID - 1):0])
    ,.a_wlast(split8_merge10_wlast)
    ,.a_wready(split8_merge10_wready)
    ,.a_wstrb(split8_merge10_wstrb[(WSTRB - 1):0])
    ,.a_wvalid(split8_merge10_wvalid)

    ,.b_araddr(split9_merge10_araddr[31:0])
    ,.b_arburst(split9_merge10_arburst[1:0])
    ,.b_arextras(split9_merge10_arextras[(EXTRAS - 1):0])
    ,.b_arid(split9_merge10_arid[(IDWID - 1):0])
    ,.b_arlen(split9_merge10_arlen[7:0])
    ,.b_arready(split9_merge10_arready)
    ,.b_arvalid(split9_merge10_arvalid)
    ,.b_awaddr(split9_merge10_awaddr[31:0])
    ,.b_awburst(split9_merge10_awburst[1:0])
    ,.b_awextras(split9_merge10_awextras[(EXTRAS - 1):0])
    ,.b_awid(split9_merge10_awid[(IDWID - 1):0])
    ,.b_awlen(split9_merge10_awlen[7:0])
    ,.b_awready(split9_merge10_awready)
    ,.b_awvalid(split9_merge10_awvalid)
    ,.b_bid(split9_merge10_bid[(IDWID - 1):0])
    ,.b_bready(split9_merge10_bready)
    ,.b_bresp(split9_merge10_bresp[1:0])
    ,.b_bvalid(split9_merge10_bvalid)
    ,.b_rdata(split9_merge10_rdata[(DWID - 1):0])
    ,.b_rid(split9_merge10_rid[(IDWID - 1):0])
    ,.b_rlast(split9_merge10_rlast)
    ,.b_rready(split9_merge10_rready)
    ,.b_rresp(split9_merge10_rresp[1:0])
    ,.b_rvalid(split9_merge10_rvalid)
    ,.b_wdata(split9_merge10_wdata[(DWID - 1):0])
    ,.b_wlast(split9_merge10_wlast)
    ,.b_wready(split9_merge10_wready)
    ,.b_wstrb(split9_merge10_wstrb[(WSTRB - 1):0])
    ,.b_wvalid(split9_merge10_wvalid)

    ,.c_araddr(split10_merge10_araddr[31:0])
    ,.c_arburst(split10_merge10_arburst[1:0])
    ,.c_arextras(split10_merge10_arextras[(EXTRAS - 1):0])
    ,.c_arid(split10_merge10_arid[(IDWID - 1):0])
    ,.c_arlen(split10_merge10_arlen[7:0])
    ,.c_arready(split10_merge10_arready)
    ,.c_arvalid(split10_merge10_arvalid)
    ,.c_awaddr(split10_merge10_awaddr[31:0])
    ,.c_awburst(split10_merge10_awburst[1:0])
    ,.c_awextras(split10_merge10_awextras[(EXTRAS - 1):0])
    ,.c_awid(split10_merge10_awid[(IDWID - 1):0])
    ,.c_awlen(split10_merge10_awlen[7:0])
    ,.c_awready(split10_merge10_awready)
    ,.c_awvalid(split10_merge10_awvalid)
    ,.c_bid(split10_merge10_bid[(IDWID - 1):0])
    ,.c_bready(split10_merge10_bready)
    ,.c_bresp(split10_merge10_bresp[1:0])
    ,.c_bvalid(split10_merge10_bvalid)
    ,.c_rdata(split10_merge10_rdata[(DWID - 1):0])
    ,.c_rid(split10_merge10_rid[(IDWID - 1):0])
    ,.c_rlast(split10_merge10_rlast)
    ,.c_rready(split10_merge10_rready)
    ,.c_rresp(split10_merge10_rresp[1:0])
    ,.c_rvalid(split10_merge10_rvalid)
    ,.c_wdata(split10_merge10_wdata[(DWID - 1):0])
    ,.c_wlast(split10_merge10_wlast)
    ,.c_wready(split10_merge10_wready)
    ,.c_wstrb(split10_merge10_wstrb[(WSTRB - 1):0])
    ,.c_wvalid(split10_merge10_wvalid)

    ,.d_araddr(split11_merge10_araddr[31:0])
    ,.d_arburst(split11_merge10_arburst[1:0])
    ,.d_arextras(split11_merge10_arextras[(EXTRAS - 1):0])
    ,.d_arid(split11_merge10_arid[(IDWID - 1):0])
    ,.d_arlen(split11_merge10_arlen[7:0])
    ,.d_arready(split11_merge10_arready)
    ,.d_arvalid(split11_merge10_arvalid)
    ,.d_awaddr(split11_merge10_awaddr[31:0])
    ,.d_awburst(split11_merge10_awburst[1:0])
    ,.d_awextras(split11_merge10_awextras[(EXTRAS - 1):0])
    ,.d_awid(split11_merge10_awid[(IDWID - 1):0])
    ,.d_awlen(split11_merge10_awlen[7:0])
    ,.d_awready(split11_merge10_awready)
    ,.d_awvalid(split11_merge10_awvalid)
    ,.d_bid(split11_merge10_bid[(IDWID - 1):0])
    ,.d_bready(split11_merge10_bready)
    ,.d_bresp(split11_merge10_bresp[1:0])
    ,.d_bvalid(split11_merge10_bvalid)
    ,.d_rdata(split11_merge10_rdata[(DWID - 1):0])
    ,.d_rid(split11_merge10_rid[(IDWID - 1):0])
    ,.d_rlast(split11_merge10_rlast)
    ,.d_rready(split11_merge10_rready)
    ,.d_rresp(split11_merge10_rresp[1:0])
    ,.d_rvalid(split11_merge10_rvalid)
    ,.d_wdata(split11_merge10_wdata[(DWID - 1):0])
    ,.d_wlast(split11_merge10_wlast)
    ,.d_wready(split11_merge10_wready)
    ,.d_wstrb(split11_merge10_wstrb[(WSTRB - 1):0])
    ,.d_wvalid(split11_merge10_wvalid)
);


wire [IDWID-1:0] merge11_split111_arid ;
wire [31:0] merge11_split111_araddr ;
wire [7:0] merge11_split111_arlen ;
wire [EXTRAS-1:0] merge11_split111_arextras ;
wire [1:0] merge11_split111_arburst ;
wire merge11_split111_arvalid ;
wire merge11_split111_arready ;
wire [IDWID-1:0] merge11_split111_rid ;
wire [DWID-1:0] merge11_split111_rdata ;
wire [1:0] merge11_split111_rresp ;
wire merge11_split111_rlast ;
wire merge11_split111_rvalid ;
wire merge11_split111_rready ;

wire [IDWID-1:0] merge11_split111_awid ;
wire [31:0] merge11_split111_awaddr ;
wire [7:0] merge11_split111_awlen ;
wire [EXTRAS-1:0] merge11_split111_awextras ;
wire [1:0] merge11_split111_awburst ;
wire merge11_split111_awvalid ;
wire merge11_split111_awready ;
wire [DWID-1:0] merge11_split111_wdata ;
wire [WSTRB-1:0] merge11_split111_wstrb ;
wire merge11_split111_wlast ;
wire merge11_split111_wvalid ;
wire merge11_split111_wready ;
wire [IDWID-1:0] merge11_split111_bid ;
wire [1:0] merge11_split111_bresp ;
wire merge11_split111_bvalid ;
wire merge11_split111_bready ;


wire [IDWID-1:0] split9_merge11_arid ;
wire [31:0] split9_merge11_araddr ;
wire [7:0] split9_merge11_arlen ;
wire [EXTRAS-1:0] split9_merge11_arextras ;
wire [1:0] split9_merge11_arburst ;
wire split9_merge11_arvalid ;
wire split9_merge11_arready ;
wire [IDWID-1:0] split9_merge11_rid ;
wire [DWID-1:0] split9_merge11_rdata ;
wire [1:0] split9_merge11_rresp ;
wire split9_merge11_rlast ;
wire split9_merge11_rvalid ;
wire split9_merge11_rready ;

wire [IDWID-1:0] split9_merge11_awid ;
wire [31:0] split9_merge11_awaddr ;
wire [7:0] split9_merge11_awlen ;
wire [EXTRAS-1:0] split9_merge11_awextras ;
wire [1:0] split9_merge11_awburst ;
wire split9_merge11_awvalid ;
wire split9_merge11_awready ;
wire [DWID-1:0] split9_merge11_wdata ;
wire [WSTRB-1:0] split9_merge11_wstrb ;
wire split9_merge11_wlast ;
wire split9_merge11_wvalid ;
wire split9_merge11_wready ;
wire [IDWID-1:0] split9_merge11_bid ;
wire [1:0] split9_merge11_bresp ;
wire split9_merge11_bvalid ;
wire split9_merge11_bready ;


wire [IDWID-1:0] split10_merge11_arid ;
wire [31:0] split10_merge11_araddr ;
wire [7:0] split10_merge11_arlen ;
wire [EXTRAS-1:0] split10_merge11_arextras ;
wire [1:0] split10_merge11_arburst ;
wire split10_merge11_arvalid ;
wire split10_merge11_arready ;
wire [IDWID-1:0] split10_merge11_rid ;
wire [DWID-1:0] split10_merge11_rdata ;
wire [1:0] split10_merge11_rresp ;
wire split10_merge11_rlast ;
wire split10_merge11_rvalid ;
wire split10_merge11_rready ;

wire [IDWID-1:0] split10_merge11_awid ;
wire [31:0] split10_merge11_awaddr ;
wire [7:0] split10_merge11_awlen ;
wire [EXTRAS-1:0] split10_merge11_awextras ;
wire [1:0] split10_merge11_awburst ;
wire split10_merge11_awvalid ;
wire split10_merge11_awready ;
wire [DWID-1:0] split10_merge11_wdata ;
wire [WSTRB-1:0] split10_merge11_wstrb ;
wire split10_merge11_wlast ;
wire split10_merge11_wvalid ;
wire split10_merge11_wready ;
wire [IDWID-1:0] split10_merge11_bid ;
wire [1:0] split10_merge11_bresp ;
wire split10_merge11_bvalid ;
wire split10_merge11_bready ;


wire [IDWID-1:0] split11_merge11_arid ;
wire [31:0] split11_merge11_araddr ;
wire [7:0] split11_merge11_arlen ;
wire [EXTRAS-1:0] split11_merge11_arextras ;
wire [1:0] split11_merge11_arburst ;
wire split11_merge11_arvalid ;
wire split11_merge11_arready ;
wire [IDWID-1:0] split11_merge11_rid ;
wire [DWID-1:0] split11_merge11_rdata ;
wire [1:0] split11_merge11_rresp ;
wire split11_merge11_rlast ;
wire split11_merge11_rvalid ;
wire split11_merge11_rready ;

wire [IDWID-1:0] split11_merge11_awid ;
wire [31:0] split11_merge11_awaddr ;
wire [7:0] split11_merge11_awlen ;
wire [EXTRAS-1:0] split11_merge11_awextras ;
wire [1:0] split11_merge11_awburst ;
wire split11_merge11_awvalid ;
wire split11_merge11_awready ;
wire [DWID-1:0] split11_merge11_wdata ;
wire [WSTRB-1:0] split11_merge11_wstrb ;
wire split11_merge11_wlast ;
wire split11_merge11_wvalid ;
wire split11_merge11_wready ;
wire [IDWID-1:0] split11_merge11_bid ;
wire [1:0] split11_merge11_bresp ;
wire split11_merge11_bvalid ;
wire split11_merge11_bready ;


axi_4_merger merge11 (
     .clk(clk),.rst_n(rst_n)
    ,.araddr(merge11_split111_araddr[31:0])
    ,.arburst(merge11_split111_arburst[1:0])
    ,.arextras(merge11_split111_arextras[(EXTRAS - 1):0])
    ,.arid(merge11_split111_arid[(IDWID - 1):0])
    ,.arlen(merge11_split111_arlen[7:0])
    ,.arready(merge11_split111_arready)
    ,.arvalid(merge11_split111_arvalid)
    ,.awaddr(merge11_split111_awaddr[31:0])
    ,.awburst(merge11_split111_awburst[1:0])
    ,.awextras(merge11_split111_awextras[(EXTRAS - 1):0])
    ,.awid(merge11_split111_awid[3:0])
    ,.awlen(merge11_split111_awlen[7:0])
    ,.awready(merge11_split111_awready)
    ,.awvalid(merge11_split111_awvalid)
    ,.bid(merge11_split111_bid[(IDWID - 1):0])
    ,.bready(merge11_split111_bready)
    ,.bresp(merge11_split111_bresp[1:0])
    ,.bvalid(merge11_split111_bvalid)
    ,.rid(merge11_split111_rid[(IDWID - 1):0])
    ,.rlast(merge11_split111_rlast)
    ,.rready(merge11_split111_rready)
    ,.rresp(merge11_split111_rresp[1:0])
    ,.rvalid(merge11_split111_rvalid)
    ,.rdata(merge11_split111_rdata[(DWID - 1):0])
    ,.wdata(merge11_split111_wdata[(DWID - 1):0])
    ,.wlast(merge11_split111_wlast)
    ,.wready(merge11_split111_wready)
    ,.wstrb(merge11_split111_wstrb[(WSTRB - 1):0])
    ,.wvalid(merge11_split111_wvalid)


    ,.a_araddr(split8_merge11_araddr[31:0])
    ,.a_arburst(split8_merge11_arburst[1:0])
    ,.a_arextras(split8_merge11_arextras[(EXTRAS - 1):0])
    ,.a_arid(split8_merge11_arid[(IDWID - 1):0])
    ,.a_arlen(split8_merge11_arlen[7:0])
    ,.a_arready(split8_merge11_arready)
    ,.a_arvalid(split8_merge11_arvalid)
    ,.a_awaddr(split8_merge11_awaddr[31:0])
    ,.a_awburst(split8_merge11_awburst[1:0])
    ,.a_awextras(split8_merge11_awextras[(EXTRAS - 1):0])
    ,.a_awid(split8_merge11_awid[(IDWID - 1):0])
    ,.a_awlen(split8_merge11_awlen[7:0])
    ,.a_awready(split8_merge11_awready)
    ,.a_awvalid(split8_merge11_awvalid)
    ,.a_bid(split8_merge11_bid[(IDWID - 1):0])
    ,.a_bready(split8_merge11_bready)
    ,.a_bresp(split8_merge11_bresp[1:0])
    ,.a_bvalid(split8_merge11_bvalid)
    ,.a_rdata(split8_merge11_rdata[(DWID - 1):0])
    ,.a_rid(split8_merge11_rid[(IDWID - 1):0])
    ,.a_rlast(split8_merge11_rlast)
    ,.a_rready(split8_merge11_rready)
    ,.a_rresp(split8_merge11_rresp[1:0])
    ,.a_rvalid(split8_merge11_rvalid)
    ,.a_wdata(split8_merge11_wdata[(DWID - 1):0])
    ,.a_wlast(split8_merge11_wlast)
    ,.a_wready(split8_merge11_wready)
    ,.a_wstrb(split8_merge11_wstrb[(WSTRB - 1):0])
    ,.a_wvalid(split8_merge11_wvalid)

    ,.b_araddr(split9_merge11_araddr[31:0])
    ,.b_arburst(split9_merge11_arburst[1:0])
    ,.b_arextras(split9_merge11_arextras[(EXTRAS - 1):0])
    ,.b_arid(split9_merge11_arid[(IDWID - 1):0])
    ,.b_arlen(split9_merge11_arlen[7:0])
    ,.b_arready(split9_merge11_arready)
    ,.b_arvalid(split9_merge11_arvalid)
    ,.b_awaddr(split9_merge11_awaddr[31:0])
    ,.b_awburst(split9_merge11_awburst[1:0])
    ,.b_awextras(split9_merge11_awextras[(EXTRAS - 1):0])
    ,.b_awid(split9_merge11_awid[(IDWID - 1):0])
    ,.b_awlen(split9_merge11_awlen[7:0])
    ,.b_awready(split9_merge11_awready)
    ,.b_awvalid(split9_merge11_awvalid)
    ,.b_bid(split9_merge11_bid[(IDWID - 1):0])
    ,.b_bready(split9_merge11_bready)
    ,.b_bresp(split9_merge11_bresp[1:0])
    ,.b_bvalid(split9_merge11_bvalid)
    ,.b_rdata(split9_merge11_rdata[(DWID - 1):0])
    ,.b_rid(split9_merge11_rid[(IDWID - 1):0])
    ,.b_rlast(split9_merge11_rlast)
    ,.b_rready(split9_merge11_rready)
    ,.b_rresp(split9_merge11_rresp[1:0])
    ,.b_rvalid(split9_merge11_rvalid)
    ,.b_wdata(split9_merge11_wdata[(DWID - 1):0])
    ,.b_wlast(split9_merge11_wlast)
    ,.b_wready(split9_merge11_wready)
    ,.b_wstrb(split9_merge11_wstrb[(WSTRB - 1):0])
    ,.b_wvalid(split9_merge11_wvalid)

    ,.c_araddr(split10_merge11_araddr[31:0])
    ,.c_arburst(split10_merge11_arburst[1:0])
    ,.c_arextras(split10_merge11_arextras[(EXTRAS - 1):0])
    ,.c_arid(split10_merge11_arid[(IDWID - 1):0])
    ,.c_arlen(split10_merge11_arlen[7:0])
    ,.c_arready(split10_merge11_arready)
    ,.c_arvalid(split10_merge11_arvalid)
    ,.c_awaddr(split10_merge11_awaddr[31:0])
    ,.c_awburst(split10_merge11_awburst[1:0])
    ,.c_awextras(split10_merge11_awextras[(EXTRAS - 1):0])
    ,.c_awid(split10_merge11_awid[(IDWID - 1):0])
    ,.c_awlen(split10_merge11_awlen[7:0])
    ,.c_awready(split10_merge11_awready)
    ,.c_awvalid(split10_merge11_awvalid)
    ,.c_bid(split10_merge11_bid[(IDWID - 1):0])
    ,.c_bready(split10_merge11_bready)
    ,.c_bresp(split10_merge11_bresp[1:0])
    ,.c_bvalid(split10_merge11_bvalid)
    ,.c_rdata(split10_merge11_rdata[(DWID - 1):0])
    ,.c_rid(split10_merge11_rid[(IDWID - 1):0])
    ,.c_rlast(split10_merge11_rlast)
    ,.c_rready(split10_merge11_rready)
    ,.c_rresp(split10_merge11_rresp[1:0])
    ,.c_rvalid(split10_merge11_rvalid)
    ,.c_wdata(split10_merge11_wdata[(DWID - 1):0])
    ,.c_wlast(split10_merge11_wlast)
    ,.c_wready(split10_merge11_wready)
    ,.c_wstrb(split10_merge11_wstrb[(WSTRB - 1):0])
    ,.c_wvalid(split10_merge11_wvalid)

    ,.d_araddr(split11_merge11_araddr[31:0])
    ,.d_arburst(split11_merge11_arburst[1:0])
    ,.d_arextras(split11_merge11_arextras[(EXTRAS - 1):0])
    ,.d_arid(split11_merge11_arid[(IDWID - 1):0])
    ,.d_arlen(split11_merge11_arlen[7:0])
    ,.d_arready(split11_merge11_arready)
    ,.d_arvalid(split11_merge11_arvalid)
    ,.d_awaddr(split11_merge11_awaddr[31:0])
    ,.d_awburst(split11_merge11_awburst[1:0])
    ,.d_awextras(split11_merge11_awextras[(EXTRAS - 1):0])
    ,.d_awid(split11_merge11_awid[(IDWID - 1):0])
    ,.d_awlen(split11_merge11_awlen[7:0])
    ,.d_awready(split11_merge11_awready)
    ,.d_awvalid(split11_merge11_awvalid)
    ,.d_bid(split11_merge11_bid[(IDWID - 1):0])
    ,.d_bready(split11_merge11_bready)
    ,.d_bresp(split11_merge11_bresp[1:0])
    ,.d_bvalid(split11_merge11_bvalid)
    ,.d_rdata(split11_merge11_rdata[(DWID - 1):0])
    ,.d_rid(split11_merge11_rid[(IDWID - 1):0])
    ,.d_rlast(split11_merge11_rlast)
    ,.d_rready(split11_merge11_rready)
    ,.d_rresp(split11_merge11_rresp[1:0])
    ,.d_rvalid(split11_merge11_rvalid)
    ,.d_wdata(split11_merge11_wdata[(DWID - 1):0])
    ,.d_wlast(split11_merge11_wlast)
    ,.d_wready(split11_merge11_wready)
    ,.d_wstrb(split11_merge11_wstrb[(WSTRB - 1):0])
    ,.d_wvalid(split11_merge11_wvalid)
);


axi_4_splitter split9 (
     .clk(clk) ,.rst_n(rst_n)

    ,.araddr(mst9_araddr[31:0])
    ,.arburst(mst9_arburst[1:0])
    ,.arextras(mst9_arextras[(EXTRAS - 1):0])
    ,.arid(mst9_arid[(IDWID - 1):0])
    ,.arlen(mst9_arlen[7:0])
    ,.arready(mst9_arready)
    ,.arvalid(mst9_arvalid)
    ,.awaddr(mst9_awaddr[31:0])
    ,.awburst(mst9_awburst[1:0])
    ,.awextras(mst9_awextras[(EXTRAS - 1):0])
    ,.awid(mst9_awid[3:0])
    ,.awlen(mst9_awlen[7:0])
    ,.awready(mst9_awready)
    ,.awvalid(mst9_awvalid)
    ,.bid(mst9_bid[(IDWID - 1):0])
    ,.bready(mst9_bready)
    ,.bresp(mst9_bresp[1:0])
    ,.bvalid(mst9_bvalid)
    ,.rdata(mst9_rdata[(DWID - 1):0])
    ,.rid(mst9_rid[(IDWID - 1):0])
    ,.rlast(mst9_rlast)
    ,.rready(mst9_rready)
    ,.rresp(mst9_rresp[1:0])
    ,.rvalid(mst9_rvalid)
    ,.wdata(mst9_wdata[(DWID - 1):0])
    ,.wlast(mst9_wlast)
    ,.wready(mst9_wready)
    ,.wstrb(mst9_wstrb[(WSTRB - 1):0])
    ,.wvalid(mst9_wvalid)

    ,.a_araddr(split9_merge8_araddr[31:0])
    ,.a_arburst(split9_merge8_arburst[1:0])
    ,.a_arextras(split9_merge8_arextras[(EXTRAS - 1):0])
    ,.a_arid(split9_merge8_arid[(IDWID - 1):0])
    ,.a_arlen(split9_merge8_arlen[7:0])
    ,.a_arready(split9_merge8_arready)
    ,.a_arvalid(split9_merge8_arvalid)
    ,.a_awaddr(split9_merge8_awaddr[31:0])
    ,.a_awburst(split9_merge8_awburst[1:0])
    ,.a_awextras(split9_merge8_awextras[(EXTRAS - 1):0])
    ,.a_awid(split9_merge8_awid[(IDWID - 1):0])
    ,.a_awlen(split9_merge8_awlen[7:0])
    ,.a_awready(split9_merge8_awready)
    ,.a_awvalid(split9_merge8_awvalid)
    ,.a_bid(split9_merge8_bid[(IDWID - 1):0])
    ,.a_bready(split9_merge8_bready)
    ,.a_bresp(split9_merge8_bresp[1:0])
    ,.a_bvalid(split9_merge8_bvalid)
    ,.a_rdata(split9_merge8_rdata[(DWID - 1):0])
    ,.a_rid(split9_merge8_rid[(IDWID - 1):0])
    ,.a_rlast(split9_merge8_rlast)
    ,.a_rready(split9_merge8_rready)
    ,.a_rresp(split9_merge8_rresp[1:0])
    ,.a_rvalid(split9_merge8_rvalid)
    ,.a_wdata(split9_merge8_wdata[(DWID - 1):0])
    ,.a_wlast(split9_merge8_wlast)
    ,.a_wready(split9_merge8_wready)
    ,.a_wstrb(split9_merge8_wstrb[(WSTRB - 1):0])
    ,.a_wvalid(split9_merge8_wvalid)
    ,.b_araddr(split9_merge9_araddr[31:0])
    ,.b_arburst(split9_merge9_arburst[1:0])
    ,.b_arextras(split9_merge9_arextras[(EXTRAS - 1):0])
    ,.b_arid(split9_merge9_arid[(IDWID - 1):0])
    ,.b_arlen(split9_merge9_arlen[7:0])
    ,.b_arready(split9_merge9_arready)
    ,.b_arvalid(split9_merge9_arvalid)
    ,.b_awaddr(split9_merge9_awaddr[31:0])
    ,.b_awburst(split9_merge9_awburst[1:0])
    ,.b_awextras(split9_merge9_awextras[(EXTRAS - 1):0])
    ,.b_awid(split9_merge9_awid[(IDWID - 1):0])
    ,.b_awlen(split9_merge9_awlen[7:0])
    ,.b_awready(split9_merge9_awready)
    ,.b_awvalid(split9_merge9_awvalid)
    ,.b_bid(split9_merge9_bid[(IDWID - 1):0])
    ,.b_bready(split9_merge9_bready)
    ,.b_bresp(split9_merge9_bresp[1:0])
    ,.b_bvalid(split9_merge9_bvalid)
    ,.b_rdata(split9_merge9_rdata[(DWID - 1):0])
    ,.b_rid(split9_merge9_rid[(IDWID - 1):0])
    ,.b_rlast(split9_merge9_rlast)
    ,.b_rready(split9_merge9_rready)
    ,.b_rresp(split9_merge9_rresp[1:0])
    ,.b_rvalid(split9_merge9_rvalid)
    ,.b_wdata(split9_merge9_wdata[(DWID - 1):0])
    ,.b_wlast(split9_merge9_wlast)
    ,.b_wready(split9_merge9_wready)
    ,.b_wstrb(split9_merge9_wstrb[(WSTRB - 1):0])
    ,.b_wvalid(split9_merge9_wvalid)
    ,.c_araddr(split9_merge10_araddr[31:0])
    ,.c_arburst(split9_merge10_arburst[1:0])
    ,.c_arextras(split9_merge10_arextras[(EXTRAS - 1):0])
    ,.c_arid(split9_merge10_arid[(IDWID - 1):0])
    ,.c_arlen(split9_merge10_arlen[7:0])
    ,.c_arready(split9_merge10_arready)
    ,.c_arvalid(split9_merge10_arvalid)
    ,.c_awaddr(split9_merge10_awaddr[31:0])
    ,.c_awburst(split9_merge10_awburst[1:0])
    ,.c_awextras(split9_merge10_awextras[(EXTRAS - 1):0])
    ,.c_awid(split9_merge10_awid[(IDWID - 1):0])
    ,.c_awlen(split9_merge10_awlen[7:0])
    ,.c_awready(split9_merge10_awready)
    ,.c_awvalid(split9_merge10_awvalid)
    ,.c_bid(split9_merge10_bid[(IDWID - 1):0])
    ,.c_bready(split9_merge10_bready)
    ,.c_bresp(split9_merge10_bresp[1:0])
    ,.c_bvalid(split9_merge10_bvalid)
    ,.c_rdata(split9_merge10_rdata[(DWID - 1):0])
    ,.c_rid(split9_merge10_rid[(IDWID - 1):0])
    ,.c_rlast(split9_merge10_rlast)
    ,.c_rready(split9_merge10_rready)
    ,.c_rresp(split9_merge10_rresp[1:0])
    ,.c_rvalid(split9_merge10_rvalid)
    ,.c_wdata(split9_merge10_wdata[(DWID - 1):0])
    ,.c_wlast(split9_merge10_wlast)
    ,.c_wready(split9_merge10_wready)
    ,.c_wstrb(split9_merge10_wstrb[(WSTRB - 1):0])
    ,.c_wvalid(split9_merge10_wvalid)
    ,.d_araddr(split9_merge11_araddr[31:0])
    ,.d_arburst(split9_merge11_arburst[1:0])
    ,.d_arextras(split9_merge11_arextras[(EXTRAS - 1):0])
    ,.d_arid(split9_merge11_arid[(IDWID - 1):0])
    ,.d_arlen(split9_merge11_arlen[7:0])
    ,.d_arready(split9_merge11_arready)
    ,.d_arvalid(split9_merge11_arvalid)
    ,.d_awaddr(split9_merge11_awaddr[31:0])
    ,.d_awburst(split9_merge11_awburst[1:0])
    ,.d_awextras(split9_merge11_awextras[(EXTRAS - 1):0])
    ,.d_awid(split9_merge11_awid[(IDWID - 1):0])
    ,.d_awlen(split9_merge11_awlen[7:0])
    ,.d_awready(split9_merge11_awready)
    ,.d_awvalid(split9_merge11_awvalid)
    ,.d_bid(split9_merge11_bid[(IDWID - 1):0])
    ,.d_bready(split9_merge11_bready)
    ,.d_bresp(split9_merge11_bresp[1:0])
    ,.d_bvalid(split9_merge11_bvalid)
    ,.d_rdata(split9_merge11_rdata[(DWID - 1):0])
    ,.d_rid(split9_merge11_rid[(IDWID - 1):0])
    ,.d_rlast(split9_merge11_rlast)
    ,.d_rready(split9_merge11_rready)
    ,.d_rresp(split9_merge11_rresp[1:0])
    ,.d_rvalid(split9_merge11_rvalid)
    ,.d_wdata(split9_merge11_wdata[(DWID - 1):0])
    ,.d_wlast(split9_merge11_wlast)
    ,.d_wready(split9_merge11_wready)
    ,.d_wstrb(split9_merge11_wstrb[(WSTRB - 1):0])
    ,.d_wvalid(split9_merge11_wvalid)

);

axi_4_splitter split10 (
     .clk(clk) ,.rst_n(rst_n)

    ,.araddr(mst10_araddr[31:0])
    ,.arburst(mst10_arburst[1:0])
    ,.arextras(mst10_arextras[(EXTRAS - 1):0])
    ,.arid(mst10_arid[(IDWID - 1):0])
    ,.arlen(mst10_arlen[7:0])
    ,.arready(mst10_arready)
    ,.arvalid(mst10_arvalid)
    ,.awaddr(mst10_awaddr[31:0])
    ,.awburst(mst10_awburst[1:0])
    ,.awextras(mst10_awextras[(EXTRAS - 1):0])
    ,.awid(mst10_awid[3:0])
    ,.awlen(mst10_awlen[7:0])
    ,.awready(mst10_awready)
    ,.awvalid(mst10_awvalid)
    ,.bid(mst10_bid[(IDWID - 1):0])
    ,.bready(mst10_bready)
    ,.bresp(mst10_bresp[1:0])
    ,.bvalid(mst10_bvalid)
    ,.rdata(mst10_rdata[(DWID - 1):0])
    ,.rid(mst10_rid[(IDWID - 1):0])
    ,.rlast(mst10_rlast)
    ,.rready(mst10_rready)
    ,.rresp(mst10_rresp[1:0])
    ,.rvalid(mst10_rvalid)
    ,.wdata(mst10_wdata[(DWID - 1):0])
    ,.wlast(mst10_wlast)
    ,.wready(mst10_wready)
    ,.wstrb(mst10_wstrb[(WSTRB - 1):0])
    ,.wvalid(mst10_wvalid)

    ,.a_araddr(split10_merge8_araddr[31:0])
    ,.a_arburst(split10_merge8_arburst[1:0])
    ,.a_arextras(split10_merge8_arextras[(EXTRAS - 1):0])
    ,.a_arid(split10_merge8_arid[(IDWID - 1):0])
    ,.a_arlen(split10_merge8_arlen[7:0])
    ,.a_arready(split10_merge8_arready)
    ,.a_arvalid(split10_merge8_arvalid)
    ,.a_awaddr(split10_merge8_awaddr[31:0])
    ,.a_awburst(split10_merge8_awburst[1:0])
    ,.a_awextras(split10_merge8_awextras[(EXTRAS - 1):0])
    ,.a_awid(split10_merge8_awid[(IDWID - 1):0])
    ,.a_awlen(split10_merge8_awlen[7:0])
    ,.a_awready(split10_merge8_awready)
    ,.a_awvalid(split10_merge8_awvalid)
    ,.a_bid(split10_merge8_bid[(IDWID - 1):0])
    ,.a_bready(split10_merge8_bready)
    ,.a_bresp(split10_merge8_bresp[1:0])
    ,.a_bvalid(split10_merge8_bvalid)
    ,.a_rdata(split10_merge8_rdata[(DWID - 1):0])
    ,.a_rid(split10_merge8_rid[(IDWID - 1):0])
    ,.a_rlast(split10_merge8_rlast)
    ,.a_rready(split10_merge8_rready)
    ,.a_rresp(split10_merge8_rresp[1:0])
    ,.a_rvalid(split10_merge8_rvalid)
    ,.a_wdata(split10_merge8_wdata[(DWID - 1):0])
    ,.a_wlast(split10_merge8_wlast)
    ,.a_wready(split10_merge8_wready)
    ,.a_wstrb(split10_merge8_wstrb[(WSTRB - 1):0])
    ,.a_wvalid(split10_merge8_wvalid)
    ,.b_araddr(split10_merge9_araddr[31:0])
    ,.b_arburst(split10_merge9_arburst[1:0])
    ,.b_arextras(split10_merge9_arextras[(EXTRAS - 1):0])
    ,.b_arid(split10_merge9_arid[(IDWID - 1):0])
    ,.b_arlen(split10_merge9_arlen[7:0])
    ,.b_arready(split10_merge9_arready)
    ,.b_arvalid(split10_merge9_arvalid)
    ,.b_awaddr(split10_merge9_awaddr[31:0])
    ,.b_awburst(split10_merge9_awburst[1:0])
    ,.b_awextras(split10_merge9_awextras[(EXTRAS - 1):0])
    ,.b_awid(split10_merge9_awid[(IDWID - 1):0])
    ,.b_awlen(split10_merge9_awlen[7:0])
    ,.b_awready(split10_merge9_awready)
    ,.b_awvalid(split10_merge9_awvalid)
    ,.b_bid(split10_merge9_bid[(IDWID - 1):0])
    ,.b_bready(split10_merge9_bready)
    ,.b_bresp(split10_merge9_bresp[1:0])
    ,.b_bvalid(split10_merge9_bvalid)
    ,.b_rdata(split10_merge9_rdata[(DWID - 1):0])
    ,.b_rid(split10_merge9_rid[(IDWID - 1):0])
    ,.b_rlast(split10_merge9_rlast)
    ,.b_rready(split10_merge9_rready)
    ,.b_rresp(split10_merge9_rresp[1:0])
    ,.b_rvalid(split10_merge9_rvalid)
    ,.b_wdata(split10_merge9_wdata[(DWID - 1):0])
    ,.b_wlast(split10_merge9_wlast)
    ,.b_wready(split10_merge9_wready)
    ,.b_wstrb(split10_merge9_wstrb[(WSTRB - 1):0])
    ,.b_wvalid(split10_merge9_wvalid)
    ,.c_araddr(split10_merge10_araddr[31:0])
    ,.c_arburst(split10_merge10_arburst[1:0])
    ,.c_arextras(split10_merge10_arextras[(EXTRAS - 1):0])
    ,.c_arid(split10_merge10_arid[(IDWID - 1):0])
    ,.c_arlen(split10_merge10_arlen[7:0])
    ,.c_arready(split10_merge10_arready)
    ,.c_arvalid(split10_merge10_arvalid)
    ,.c_awaddr(split10_merge10_awaddr[31:0])
    ,.c_awburst(split10_merge10_awburst[1:0])
    ,.c_awextras(split10_merge10_awextras[(EXTRAS - 1):0])
    ,.c_awid(split10_merge10_awid[(IDWID - 1):0])
    ,.c_awlen(split10_merge10_awlen[7:0])
    ,.c_awready(split10_merge10_awready)
    ,.c_awvalid(split10_merge10_awvalid)
    ,.c_bid(split10_merge10_bid[(IDWID - 1):0])
    ,.c_bready(split10_merge10_bready)
    ,.c_bresp(split10_merge10_bresp[1:0])
    ,.c_bvalid(split10_merge10_bvalid)
    ,.c_rdata(split10_merge10_rdata[(DWID - 1):0])
    ,.c_rid(split10_merge10_rid[(IDWID - 1):0])
    ,.c_rlast(split10_merge10_rlast)
    ,.c_rready(split10_merge10_rready)
    ,.c_rresp(split10_merge10_rresp[1:0])
    ,.c_rvalid(split10_merge10_rvalid)
    ,.c_wdata(split10_merge10_wdata[(DWID - 1):0])
    ,.c_wlast(split10_merge10_wlast)
    ,.c_wready(split10_merge10_wready)
    ,.c_wstrb(split10_merge10_wstrb[(WSTRB - 1):0])
    ,.c_wvalid(split10_merge10_wvalid)
    ,.d_araddr(split10_merge11_araddr[31:0])
    ,.d_arburst(split10_merge11_arburst[1:0])
    ,.d_arextras(split10_merge11_arextras[(EXTRAS - 1):0])
    ,.d_arid(split10_merge11_arid[(IDWID - 1):0])
    ,.d_arlen(split10_merge11_arlen[7:0])
    ,.d_arready(split10_merge11_arready)
    ,.d_arvalid(split10_merge11_arvalid)
    ,.d_awaddr(split10_merge11_awaddr[31:0])
    ,.d_awburst(split10_merge11_awburst[1:0])
    ,.d_awextras(split10_merge11_awextras[(EXTRAS - 1):0])
    ,.d_awid(split10_merge11_awid[(IDWID - 1):0])
    ,.d_awlen(split10_merge11_awlen[7:0])
    ,.d_awready(split10_merge11_awready)
    ,.d_awvalid(split10_merge11_awvalid)
    ,.d_bid(split10_merge11_bid[(IDWID - 1):0])
    ,.d_bready(split10_merge11_bready)
    ,.d_bresp(split10_merge11_bresp[1:0])
    ,.d_bvalid(split10_merge11_bvalid)
    ,.d_rdata(split10_merge11_rdata[(DWID - 1):0])
    ,.d_rid(split10_merge11_rid[(IDWID - 1):0])
    ,.d_rlast(split10_merge11_rlast)
    ,.d_rready(split10_merge11_rready)
    ,.d_rresp(split10_merge11_rresp[1:0])
    ,.d_rvalid(split10_merge11_rvalid)
    ,.d_wdata(split10_merge11_wdata[(DWID - 1):0])
    ,.d_wlast(split10_merge11_wlast)
    ,.d_wready(split10_merge11_wready)
    ,.d_wstrb(split10_merge11_wstrb[(WSTRB - 1):0])
    ,.d_wvalid(split10_merge11_wvalid)

);

axi_4_splitter split11 (
     .clk(clk) ,.rst_n(rst_n)

    ,.araddr(mst11_araddr[31:0])
    ,.arburst(mst11_arburst[1:0])
    ,.arextras(mst11_arextras[(EXTRAS - 1):0])
    ,.arid(mst11_arid[(IDWID - 1):0])
    ,.arlen(mst11_arlen[7:0])
    ,.arready(mst11_arready)
    ,.arvalid(mst11_arvalid)
    ,.awaddr(mst11_awaddr[31:0])
    ,.awburst(mst11_awburst[1:0])
    ,.awextras(mst11_awextras[(EXTRAS - 1):0])
    ,.awid(mst11_awid[3:0])
    ,.awlen(mst11_awlen[7:0])
    ,.awready(mst11_awready)
    ,.awvalid(mst11_awvalid)
    ,.bid(mst11_bid[(IDWID - 1):0])
    ,.bready(mst11_bready)
    ,.bresp(mst11_bresp[1:0])
    ,.bvalid(mst11_bvalid)
    ,.rdata(mst11_rdata[(DWID - 1):0])
    ,.rid(mst11_rid[(IDWID - 1):0])
    ,.rlast(mst11_rlast)
    ,.rready(mst11_rready)
    ,.rresp(mst11_rresp[1:0])
    ,.rvalid(mst11_rvalid)
    ,.wdata(mst11_wdata[(DWID - 1):0])
    ,.wlast(mst11_wlast)
    ,.wready(mst11_wready)
    ,.wstrb(mst11_wstrb[(WSTRB - 1):0])
    ,.wvalid(mst11_wvalid)

    ,.a_araddr(split11_merge8_araddr[31:0])
    ,.a_arburst(split11_merge8_arburst[1:0])
    ,.a_arextras(split11_merge8_arextras[(EXTRAS - 1):0])
    ,.a_arid(split11_merge8_arid[(IDWID - 1):0])
    ,.a_arlen(split11_merge8_arlen[7:0])
    ,.a_arready(split11_merge8_arready)
    ,.a_arvalid(split11_merge8_arvalid)
    ,.a_awaddr(split11_merge8_awaddr[31:0])
    ,.a_awburst(split11_merge8_awburst[1:0])
    ,.a_awextras(split11_merge8_awextras[(EXTRAS - 1):0])
    ,.a_awid(split11_merge8_awid[(IDWID - 1):0])
    ,.a_awlen(split11_merge8_awlen[7:0])
    ,.a_awready(split11_merge8_awready)
    ,.a_awvalid(split11_merge8_awvalid)
    ,.a_bid(split11_merge8_bid[(IDWID - 1):0])
    ,.a_bready(split11_merge8_bready)
    ,.a_bresp(split11_merge8_bresp[1:0])
    ,.a_bvalid(split11_merge8_bvalid)
    ,.a_rdata(split11_merge8_rdata[(DWID - 1):0])
    ,.a_rid(split11_merge8_rid[(IDWID - 1):0])
    ,.a_rlast(split11_merge8_rlast)
    ,.a_rready(split11_merge8_rready)
    ,.a_rresp(split11_merge8_rresp[1:0])
    ,.a_rvalid(split11_merge8_rvalid)
    ,.a_wdata(split11_merge8_wdata[(DWID - 1):0])
    ,.a_wlast(split11_merge8_wlast)
    ,.a_wready(split11_merge8_wready)
    ,.a_wstrb(split11_merge8_wstrb[(WSTRB - 1):0])
    ,.a_wvalid(split11_merge8_wvalid)
    ,.b_araddr(split11_merge9_araddr[31:0])
    ,.b_arburst(split11_merge9_arburst[1:0])
    ,.b_arextras(split11_merge9_arextras[(EXTRAS - 1):0])
    ,.b_arid(split11_merge9_arid[(IDWID - 1):0])
    ,.b_arlen(split11_merge9_arlen[7:0])
    ,.b_arready(split11_merge9_arready)
    ,.b_arvalid(split11_merge9_arvalid)
    ,.b_awaddr(split11_merge9_awaddr[31:0])
    ,.b_awburst(split11_merge9_awburst[1:0])
    ,.b_awextras(split11_merge9_awextras[(EXTRAS - 1):0])
    ,.b_awid(split11_merge9_awid[(IDWID - 1):0])
    ,.b_awlen(split11_merge9_awlen[7:0])
    ,.b_awready(split11_merge9_awready)
    ,.b_awvalid(split11_merge9_awvalid)
    ,.b_bid(split11_merge9_bid[(IDWID - 1):0])
    ,.b_bready(split11_merge9_bready)
    ,.b_bresp(split11_merge9_bresp[1:0])
    ,.b_bvalid(split11_merge9_bvalid)
    ,.b_rdata(split11_merge9_rdata[(DWID - 1):0])
    ,.b_rid(split11_merge9_rid[(IDWID - 1):0])
    ,.b_rlast(split11_merge9_rlast)
    ,.b_rready(split11_merge9_rready)
    ,.b_rresp(split11_merge9_rresp[1:0])
    ,.b_rvalid(split11_merge9_rvalid)
    ,.b_wdata(split11_merge9_wdata[(DWID - 1):0])
    ,.b_wlast(split11_merge9_wlast)
    ,.b_wready(split11_merge9_wready)
    ,.b_wstrb(split11_merge9_wstrb[(WSTRB - 1):0])
    ,.b_wvalid(split11_merge9_wvalid)
    ,.c_araddr(split11_merge10_araddr[31:0])
    ,.c_arburst(split11_merge10_arburst[1:0])
    ,.c_arextras(split11_merge10_arextras[(EXTRAS - 1):0])
    ,.c_arid(split11_merge10_arid[(IDWID - 1):0])
    ,.c_arlen(split11_merge10_arlen[7:0])
    ,.c_arready(split11_merge10_arready)
    ,.c_arvalid(split11_merge10_arvalid)
    ,.c_awaddr(split11_merge10_awaddr[31:0])
    ,.c_awburst(split11_merge10_awburst[1:0])
    ,.c_awextras(split11_merge10_awextras[(EXTRAS - 1):0])
    ,.c_awid(split11_merge10_awid[(IDWID - 1):0])
    ,.c_awlen(split11_merge10_awlen[7:0])
    ,.c_awready(split11_merge10_awready)
    ,.c_awvalid(split11_merge10_awvalid)
    ,.c_bid(split11_merge10_bid[(IDWID - 1):0])
    ,.c_bready(split11_merge10_bready)
    ,.c_bresp(split11_merge10_bresp[1:0])
    ,.c_bvalid(split11_merge10_bvalid)
    ,.c_rdata(split11_merge10_rdata[(DWID - 1):0])
    ,.c_rid(split11_merge10_rid[(IDWID - 1):0])
    ,.c_rlast(split11_merge10_rlast)
    ,.c_rready(split11_merge10_rready)
    ,.c_rresp(split11_merge10_rresp[1:0])
    ,.c_rvalid(split11_merge10_rvalid)
    ,.c_wdata(split11_merge10_wdata[(DWID - 1):0])
    ,.c_wlast(split11_merge10_wlast)
    ,.c_wready(split11_merge10_wready)
    ,.c_wstrb(split11_merge10_wstrb[(WSTRB - 1):0])
    ,.c_wvalid(split11_merge10_wvalid)
    ,.d_araddr(split11_merge11_araddr[31:0])
    ,.d_arburst(split11_merge11_arburst[1:0])
    ,.d_arextras(split11_merge11_arextras[(EXTRAS - 1):0])
    ,.d_arid(split11_merge11_arid[(IDWID - 1):0])
    ,.d_arlen(split11_merge11_arlen[7:0])
    ,.d_arready(split11_merge11_arready)
    ,.d_arvalid(split11_merge11_arvalid)
    ,.d_awaddr(split11_merge11_awaddr[31:0])
    ,.d_awburst(split11_merge11_awburst[1:0])
    ,.d_awextras(split11_merge11_awextras[(EXTRAS - 1):0])
    ,.d_awid(split11_merge11_awid[(IDWID - 1):0])
    ,.d_awlen(split11_merge11_awlen[7:0])
    ,.d_awready(split11_merge11_awready)
    ,.d_awvalid(split11_merge11_awvalid)
    ,.d_bid(split11_merge11_bid[(IDWID - 1):0])
    ,.d_bready(split11_merge11_bready)
    ,.d_bresp(split11_merge11_bresp[1:0])
    ,.d_bvalid(split11_merge11_bvalid)
    ,.d_rdata(split11_merge11_rdata[(DWID - 1):0])
    ,.d_rid(split11_merge11_rid[(IDWID - 1):0])
    ,.d_rlast(split11_merge11_rlast)
    ,.d_rready(split11_merge11_rready)
    ,.d_rresp(split11_merge11_rresp[1:0])
    ,.d_rvalid(split11_merge11_rvalid)
    ,.d_wdata(split11_merge11_wdata[(DWID - 1):0])
    ,.d_wlast(split11_merge11_wlast)
    ,.d_wready(split11_merge11_wready)
    ,.d_wstrb(split11_merge11_wstrb[(WSTRB - 1):0])
    ,.d_wvalid(split11_merge11_wvalid)

);

wire [IDWID-1:0] split12_merge12_arid ;
wire [31:0] split12_merge12_araddr ;
wire [7:0] split12_merge12_arlen ;
wire [EXTRAS-1:0] split12_merge12_arextras ;
wire [1:0] split12_merge12_arburst ;
wire split12_merge12_arvalid ;
wire split12_merge12_arready ;
wire [IDWID-1:0] split12_merge12_rid ;
wire [DWID-1:0] split12_merge12_rdata ;
wire [1:0] split12_merge12_rresp ;
wire split12_merge12_rlast ;
wire split12_merge12_rvalid ;
wire split12_merge12_rready ;

wire [IDWID-1:0] split12_merge12_awid ;
wire [31:0] split12_merge12_awaddr ;
wire [7:0] split12_merge12_awlen ;
wire [EXTRAS-1:0] split12_merge12_awextras ;
wire [1:0] split12_merge12_awburst ;
wire split12_merge12_awvalid ;
wire split12_merge12_awready ;
wire [DWID-1:0] split12_merge12_wdata ;
wire [WSTRB-1:0] split12_merge12_wstrb ;
wire split12_merge12_wlast ;
wire split12_merge12_wvalid ;
wire split12_merge12_wready ;
wire [IDWID-1:0] split12_merge12_bid ;
wire [1:0] split12_merge12_bresp ;
wire split12_merge12_bvalid ;
wire split12_merge12_bready ;


wire [IDWID-1:0] split12_merge13_arid ;
wire [31:0] split12_merge13_araddr ;
wire [7:0] split12_merge13_arlen ;
wire [EXTRAS-1:0] split12_merge13_arextras ;
wire [1:0] split12_merge13_arburst ;
wire split12_merge13_arvalid ;
wire split12_merge13_arready ;
wire [IDWID-1:0] split12_merge13_rid ;
wire [DWID-1:0] split12_merge13_rdata ;
wire [1:0] split12_merge13_rresp ;
wire split12_merge13_rlast ;
wire split12_merge13_rvalid ;
wire split12_merge13_rready ;

wire [IDWID-1:0] split12_merge13_awid ;
wire [31:0] split12_merge13_awaddr ;
wire [7:0] split12_merge13_awlen ;
wire [EXTRAS-1:0] split12_merge13_awextras ;
wire [1:0] split12_merge13_awburst ;
wire split12_merge13_awvalid ;
wire split12_merge13_awready ;
wire [DWID-1:0] split12_merge13_wdata ;
wire [WSTRB-1:0] split12_merge13_wstrb ;
wire split12_merge13_wlast ;
wire split12_merge13_wvalid ;
wire split12_merge13_wready ;
wire [IDWID-1:0] split12_merge13_bid ;
wire [1:0] split12_merge13_bresp ;
wire split12_merge13_bvalid ;
wire split12_merge13_bready ;


wire [IDWID-1:0] split12_merge14_arid ;
wire [31:0] split12_merge14_araddr ;
wire [7:0] split12_merge14_arlen ;
wire [EXTRAS-1:0] split12_merge14_arextras ;
wire [1:0] split12_merge14_arburst ;
wire split12_merge14_arvalid ;
wire split12_merge14_arready ;
wire [IDWID-1:0] split12_merge14_rid ;
wire [DWID-1:0] split12_merge14_rdata ;
wire [1:0] split12_merge14_rresp ;
wire split12_merge14_rlast ;
wire split12_merge14_rvalid ;
wire split12_merge14_rready ;

wire [IDWID-1:0] split12_merge14_awid ;
wire [31:0] split12_merge14_awaddr ;
wire [7:0] split12_merge14_awlen ;
wire [EXTRAS-1:0] split12_merge14_awextras ;
wire [1:0] split12_merge14_awburst ;
wire split12_merge14_awvalid ;
wire split12_merge14_awready ;
wire [DWID-1:0] split12_merge14_wdata ;
wire [WSTRB-1:0] split12_merge14_wstrb ;
wire split12_merge14_wlast ;
wire split12_merge14_wvalid ;
wire split12_merge14_wready ;
wire [IDWID-1:0] split12_merge14_bid ;
wire [1:0] split12_merge14_bresp ;
wire split12_merge14_bvalid ;
wire split12_merge14_bready ;


wire [IDWID-1:0] split12_merge15_arid ;
wire [31:0] split12_merge15_araddr ;
wire [7:0] split12_merge15_arlen ;
wire [EXTRAS-1:0] split12_merge15_arextras ;
wire [1:0] split12_merge15_arburst ;
wire split12_merge15_arvalid ;
wire split12_merge15_arready ;
wire [IDWID-1:0] split12_merge15_rid ;
wire [DWID-1:0] split12_merge15_rdata ;
wire [1:0] split12_merge15_rresp ;
wire split12_merge15_rlast ;
wire split12_merge15_rvalid ;
wire split12_merge15_rready ;

wire [IDWID-1:0] split12_merge15_awid ;
wire [31:0] split12_merge15_awaddr ;
wire [7:0] split12_merge15_awlen ;
wire [EXTRAS-1:0] split12_merge15_awextras ;
wire [1:0] split12_merge15_awburst ;
wire split12_merge15_awvalid ;
wire split12_merge15_awready ;
wire [DWID-1:0] split12_merge15_wdata ;
wire [WSTRB-1:0] split12_merge15_wstrb ;
wire split12_merge15_wlast ;
wire split12_merge15_wvalid ;
wire split12_merge15_wready ;
wire [IDWID-1:0] split12_merge15_bid ;
wire [1:0] split12_merge15_bresp ;
wire split12_merge15_bvalid ;
wire split12_merge15_bready ;


axi_4_splitter split12 (
     .clk(clk) ,.rst_n(rst_n)

    ,.araddr(mst12_araddr[31:0])
    ,.arburst(mst12_arburst[1:0])
    ,.arextras(mst12_arextras[(EXTRAS - 1):0])
    ,.arid(mst12_arid[(IDWID - 1):0])
    ,.arlen(mst12_arlen[7:0])
    ,.arready(mst12_arready)
    ,.arvalid(mst12_arvalid)
    ,.awaddr(mst12_awaddr[31:0])
    ,.awburst(mst12_awburst[1:0])
    ,.awextras(mst12_awextras[(EXTRAS - 1):0])
    ,.awid(mst12_awid[3:0])
    ,.awlen(mst12_awlen[7:0])
    ,.awready(mst12_awready)
    ,.awvalid(mst12_awvalid)
    ,.bid(mst12_bid[(IDWID - 1):0])
    ,.bready(mst12_bready)
    ,.bresp(mst12_bresp[1:0])
    ,.bvalid(mst12_bvalid)
    ,.rdata(mst12_rdata[(DWID - 1):0])
    ,.rid(mst12_rid[(IDWID - 1):0])
    ,.rlast(mst12_rlast)
    ,.rready(mst12_rready)
    ,.rresp(mst12_rresp[1:0])
    ,.rvalid(mst12_rvalid)
    ,.wdata(mst12_wdata[(DWID - 1):0])
    ,.wlast(mst12_wlast)
    ,.wready(mst12_wready)
    ,.wstrb(mst12_wstrb[(WSTRB - 1):0])
    ,.wvalid(mst12_wvalid)

    ,.a_araddr(split12_merge12_araddr[31:0])
    ,.a_arburst(split12_merge12_arburst[1:0])
    ,.a_arextras(split12_merge12_arextras[(EXTRAS - 1):0])
    ,.a_arid(split12_merge12_arid[(IDWID - 1):0])
    ,.a_arlen(split12_merge12_arlen[7:0])
    ,.a_arready(split12_merge12_arready)
    ,.a_arvalid(split12_merge12_arvalid)
    ,.a_awaddr(split12_merge12_awaddr[31:0])
    ,.a_awburst(split12_merge12_awburst[1:0])
    ,.a_awextras(split12_merge12_awextras[(EXTRAS - 1):0])
    ,.a_awid(split12_merge12_awid[(IDWID - 1):0])
    ,.a_awlen(split12_merge12_awlen[7:0])
    ,.a_awready(split12_merge12_awready)
    ,.a_awvalid(split12_merge12_awvalid)
    ,.a_bid(split12_merge12_bid[(IDWID - 1):0])
    ,.a_bready(split12_merge12_bready)
    ,.a_bresp(split12_merge12_bresp[1:0])
    ,.a_bvalid(split12_merge12_bvalid)
    ,.a_rdata(split12_merge12_rdata[(DWID - 1):0])
    ,.a_rid(split12_merge12_rid[(IDWID - 1):0])
    ,.a_rlast(split12_merge12_rlast)
    ,.a_rready(split12_merge12_rready)
    ,.a_rresp(split12_merge12_rresp[1:0])
    ,.a_rvalid(split12_merge12_rvalid)
    ,.a_wdata(split12_merge12_wdata[(DWID - 1):0])
    ,.a_wlast(split12_merge12_wlast)
    ,.a_wready(split12_merge12_wready)
    ,.a_wstrb(split12_merge12_wstrb[(WSTRB - 1):0])
    ,.a_wvalid(split12_merge12_wvalid)
    ,.b_araddr(split12_merge13_araddr[31:0])
    ,.b_arburst(split12_merge13_arburst[1:0])
    ,.b_arextras(split12_merge13_arextras[(EXTRAS - 1):0])
    ,.b_arid(split12_merge13_arid[(IDWID - 1):0])
    ,.b_arlen(split12_merge13_arlen[7:0])
    ,.b_arready(split12_merge13_arready)
    ,.b_arvalid(split12_merge13_arvalid)
    ,.b_awaddr(split12_merge13_awaddr[31:0])
    ,.b_awburst(split12_merge13_awburst[1:0])
    ,.b_awextras(split12_merge13_awextras[(EXTRAS - 1):0])
    ,.b_awid(split12_merge13_awid[(IDWID - 1):0])
    ,.b_awlen(split12_merge13_awlen[7:0])
    ,.b_awready(split12_merge13_awready)
    ,.b_awvalid(split12_merge13_awvalid)
    ,.b_bid(split12_merge13_bid[(IDWID - 1):0])
    ,.b_bready(split12_merge13_bready)
    ,.b_bresp(split12_merge13_bresp[1:0])
    ,.b_bvalid(split12_merge13_bvalid)
    ,.b_rdata(split12_merge13_rdata[(DWID - 1):0])
    ,.b_rid(split12_merge13_rid[(IDWID - 1):0])
    ,.b_rlast(split12_merge13_rlast)
    ,.b_rready(split12_merge13_rready)
    ,.b_rresp(split12_merge13_rresp[1:0])
    ,.b_rvalid(split12_merge13_rvalid)
    ,.b_wdata(split12_merge13_wdata[(DWID - 1):0])
    ,.b_wlast(split12_merge13_wlast)
    ,.b_wready(split12_merge13_wready)
    ,.b_wstrb(split12_merge13_wstrb[(WSTRB - 1):0])
    ,.b_wvalid(split12_merge13_wvalid)
    ,.c_araddr(split12_merge14_araddr[31:0])
    ,.c_arburst(split12_merge14_arburst[1:0])
    ,.c_arextras(split12_merge14_arextras[(EXTRAS - 1):0])
    ,.c_arid(split12_merge14_arid[(IDWID - 1):0])
    ,.c_arlen(split12_merge14_arlen[7:0])
    ,.c_arready(split12_merge14_arready)
    ,.c_arvalid(split12_merge14_arvalid)
    ,.c_awaddr(split12_merge14_awaddr[31:0])
    ,.c_awburst(split12_merge14_awburst[1:0])
    ,.c_awextras(split12_merge14_awextras[(EXTRAS - 1):0])
    ,.c_awid(split12_merge14_awid[(IDWID - 1):0])
    ,.c_awlen(split12_merge14_awlen[7:0])
    ,.c_awready(split12_merge14_awready)
    ,.c_awvalid(split12_merge14_awvalid)
    ,.c_bid(split12_merge14_bid[(IDWID - 1):0])
    ,.c_bready(split12_merge14_bready)
    ,.c_bresp(split12_merge14_bresp[1:0])
    ,.c_bvalid(split12_merge14_bvalid)
    ,.c_rdata(split12_merge14_rdata[(DWID - 1):0])
    ,.c_rid(split12_merge14_rid[(IDWID - 1):0])
    ,.c_rlast(split12_merge14_rlast)
    ,.c_rready(split12_merge14_rready)
    ,.c_rresp(split12_merge14_rresp[1:0])
    ,.c_rvalid(split12_merge14_rvalid)
    ,.c_wdata(split12_merge14_wdata[(DWID - 1):0])
    ,.c_wlast(split12_merge14_wlast)
    ,.c_wready(split12_merge14_wready)
    ,.c_wstrb(split12_merge14_wstrb[(WSTRB - 1):0])
    ,.c_wvalid(split12_merge14_wvalid)
    ,.d_araddr(split12_merge15_araddr[31:0])
    ,.d_arburst(split12_merge15_arburst[1:0])
    ,.d_arextras(split12_merge15_arextras[(EXTRAS - 1):0])
    ,.d_arid(split12_merge15_arid[(IDWID - 1):0])
    ,.d_arlen(split12_merge15_arlen[7:0])
    ,.d_arready(split12_merge15_arready)
    ,.d_arvalid(split12_merge15_arvalid)
    ,.d_awaddr(split12_merge15_awaddr[31:0])
    ,.d_awburst(split12_merge15_awburst[1:0])
    ,.d_awextras(split12_merge15_awextras[(EXTRAS - 1):0])
    ,.d_awid(split12_merge15_awid[(IDWID - 1):0])
    ,.d_awlen(split12_merge15_awlen[7:0])
    ,.d_awready(split12_merge15_awready)
    ,.d_awvalid(split12_merge15_awvalid)
    ,.d_bid(split12_merge15_bid[(IDWID - 1):0])
    ,.d_bready(split12_merge15_bready)
    ,.d_bresp(split12_merge15_bresp[1:0])
    ,.d_bvalid(split12_merge15_bvalid)
    ,.d_rdata(split12_merge15_rdata[(DWID - 1):0])
    ,.d_rid(split12_merge15_rid[(IDWID - 1):0])
    ,.d_rlast(split12_merge15_rlast)
    ,.d_rready(split12_merge15_rready)
    ,.d_rresp(split12_merge15_rresp[1:0])
    ,.d_rvalid(split12_merge15_rvalid)
    ,.d_wdata(split12_merge15_wdata[(DWID - 1):0])
    ,.d_wlast(split12_merge15_wlast)
    ,.d_wready(split12_merge15_wready)
    ,.d_wstrb(split12_merge15_wstrb[(WSTRB - 1):0])
    ,.d_wvalid(split12_merge15_wvalid)

);

wire [IDWID-1:0] merge12_split112_arid ;
wire [31:0] merge12_split112_araddr ;
wire [7:0] merge12_split112_arlen ;
wire [EXTRAS-1:0] merge12_split112_arextras ;
wire [1:0] merge12_split112_arburst ;
wire merge12_split112_arvalid ;
wire merge12_split112_arready ;
wire [IDWID-1:0] merge12_split112_rid ;
wire [DWID-1:0] merge12_split112_rdata ;
wire [1:0] merge12_split112_rresp ;
wire merge12_split112_rlast ;
wire merge12_split112_rvalid ;
wire merge12_split112_rready ;

wire [IDWID-1:0] merge12_split112_awid ;
wire [31:0] merge12_split112_awaddr ;
wire [7:0] merge12_split112_awlen ;
wire [EXTRAS-1:0] merge12_split112_awextras ;
wire [1:0] merge12_split112_awburst ;
wire merge12_split112_awvalid ;
wire merge12_split112_awready ;
wire [DWID-1:0] merge12_split112_wdata ;
wire [WSTRB-1:0] merge12_split112_wstrb ;
wire merge12_split112_wlast ;
wire merge12_split112_wvalid ;
wire merge12_split112_wready ;
wire [IDWID-1:0] merge12_split112_bid ;
wire [1:0] merge12_split112_bresp ;
wire merge12_split112_bvalid ;
wire merge12_split112_bready ;


wire [IDWID-1:0] split13_merge12_arid ;
wire [31:0] split13_merge12_araddr ;
wire [7:0] split13_merge12_arlen ;
wire [EXTRAS-1:0] split13_merge12_arextras ;
wire [1:0] split13_merge12_arburst ;
wire split13_merge12_arvalid ;
wire split13_merge12_arready ;
wire [IDWID-1:0] split13_merge12_rid ;
wire [DWID-1:0] split13_merge12_rdata ;
wire [1:0] split13_merge12_rresp ;
wire split13_merge12_rlast ;
wire split13_merge12_rvalid ;
wire split13_merge12_rready ;

wire [IDWID-1:0] split13_merge12_awid ;
wire [31:0] split13_merge12_awaddr ;
wire [7:0] split13_merge12_awlen ;
wire [EXTRAS-1:0] split13_merge12_awextras ;
wire [1:0] split13_merge12_awburst ;
wire split13_merge12_awvalid ;
wire split13_merge12_awready ;
wire [DWID-1:0] split13_merge12_wdata ;
wire [WSTRB-1:0] split13_merge12_wstrb ;
wire split13_merge12_wlast ;
wire split13_merge12_wvalid ;
wire split13_merge12_wready ;
wire [IDWID-1:0] split13_merge12_bid ;
wire [1:0] split13_merge12_bresp ;
wire split13_merge12_bvalid ;
wire split13_merge12_bready ;


wire [IDWID-1:0] split14_merge12_arid ;
wire [31:0] split14_merge12_araddr ;
wire [7:0] split14_merge12_arlen ;
wire [EXTRAS-1:0] split14_merge12_arextras ;
wire [1:0] split14_merge12_arburst ;
wire split14_merge12_arvalid ;
wire split14_merge12_arready ;
wire [IDWID-1:0] split14_merge12_rid ;
wire [DWID-1:0] split14_merge12_rdata ;
wire [1:0] split14_merge12_rresp ;
wire split14_merge12_rlast ;
wire split14_merge12_rvalid ;
wire split14_merge12_rready ;

wire [IDWID-1:0] split14_merge12_awid ;
wire [31:0] split14_merge12_awaddr ;
wire [7:0] split14_merge12_awlen ;
wire [EXTRAS-1:0] split14_merge12_awextras ;
wire [1:0] split14_merge12_awburst ;
wire split14_merge12_awvalid ;
wire split14_merge12_awready ;
wire [DWID-1:0] split14_merge12_wdata ;
wire [WSTRB-1:0] split14_merge12_wstrb ;
wire split14_merge12_wlast ;
wire split14_merge12_wvalid ;
wire split14_merge12_wready ;
wire [IDWID-1:0] split14_merge12_bid ;
wire [1:0] split14_merge12_bresp ;
wire split14_merge12_bvalid ;
wire split14_merge12_bready ;


wire [IDWID-1:0] split15_merge12_arid ;
wire [31:0] split15_merge12_araddr ;
wire [7:0] split15_merge12_arlen ;
wire [EXTRAS-1:0] split15_merge12_arextras ;
wire [1:0] split15_merge12_arburst ;
wire split15_merge12_arvalid ;
wire split15_merge12_arready ;
wire [IDWID-1:0] split15_merge12_rid ;
wire [DWID-1:0] split15_merge12_rdata ;
wire [1:0] split15_merge12_rresp ;
wire split15_merge12_rlast ;
wire split15_merge12_rvalid ;
wire split15_merge12_rready ;

wire [IDWID-1:0] split15_merge12_awid ;
wire [31:0] split15_merge12_awaddr ;
wire [7:0] split15_merge12_awlen ;
wire [EXTRAS-1:0] split15_merge12_awextras ;
wire [1:0] split15_merge12_awburst ;
wire split15_merge12_awvalid ;
wire split15_merge12_awready ;
wire [DWID-1:0] split15_merge12_wdata ;
wire [WSTRB-1:0] split15_merge12_wstrb ;
wire split15_merge12_wlast ;
wire split15_merge12_wvalid ;
wire split15_merge12_wready ;
wire [IDWID-1:0] split15_merge12_bid ;
wire [1:0] split15_merge12_bresp ;
wire split15_merge12_bvalid ;
wire split15_merge12_bready ;


axi_4_merger merge12 (
     .clk(clk),.rst_n(rst_n)
    ,.araddr(merge12_split112_araddr[31:0])
    ,.arburst(merge12_split112_arburst[1:0])
    ,.arextras(merge12_split112_arextras[(EXTRAS - 1):0])
    ,.arid(merge12_split112_arid[(IDWID - 1):0])
    ,.arlen(merge12_split112_arlen[7:0])
    ,.arready(merge12_split112_arready)
    ,.arvalid(merge12_split112_arvalid)
    ,.awaddr(merge12_split112_awaddr[31:0])
    ,.awburst(merge12_split112_awburst[1:0])
    ,.awextras(merge12_split112_awextras[(EXTRAS - 1):0])
    ,.awid(merge12_split112_awid[3:0])
    ,.awlen(merge12_split112_awlen[7:0])
    ,.awready(merge12_split112_awready)
    ,.awvalid(merge12_split112_awvalid)
    ,.bid(merge12_split112_bid[(IDWID - 1):0])
    ,.bready(merge12_split112_bready)
    ,.bresp(merge12_split112_bresp[1:0])
    ,.bvalid(merge12_split112_bvalid)
    ,.rid(merge12_split112_rid[(IDWID - 1):0])
    ,.rlast(merge12_split112_rlast)
    ,.rready(merge12_split112_rready)
    ,.rresp(merge12_split112_rresp[1:0])
    ,.rvalid(merge12_split112_rvalid)
    ,.rdata(merge12_split112_rdata[(DWID - 1):0])
    ,.wdata(merge12_split112_wdata[(DWID - 1):0])
    ,.wlast(merge12_split112_wlast)
    ,.wready(merge12_split112_wready)
    ,.wstrb(merge12_split112_wstrb[(WSTRB - 1):0])
    ,.wvalid(merge12_split112_wvalid)


    ,.a_araddr(split12_merge12_araddr[31:0])
    ,.a_arburst(split12_merge12_arburst[1:0])
    ,.a_arextras(split12_merge12_arextras[(EXTRAS - 1):0])
    ,.a_arid(split12_merge12_arid[(IDWID - 1):0])
    ,.a_arlen(split12_merge12_arlen[7:0])
    ,.a_arready(split12_merge12_arready)
    ,.a_arvalid(split12_merge12_arvalid)
    ,.a_awaddr(split12_merge12_awaddr[31:0])
    ,.a_awburst(split12_merge12_awburst[1:0])
    ,.a_awextras(split12_merge12_awextras[(EXTRAS - 1):0])
    ,.a_awid(split12_merge12_awid[(IDWID - 1):0])
    ,.a_awlen(split12_merge12_awlen[7:0])
    ,.a_awready(split12_merge12_awready)
    ,.a_awvalid(split12_merge12_awvalid)
    ,.a_bid(split12_merge12_bid[(IDWID - 1):0])
    ,.a_bready(split12_merge12_bready)
    ,.a_bresp(split12_merge12_bresp[1:0])
    ,.a_bvalid(split12_merge12_bvalid)
    ,.a_rdata(split12_merge12_rdata[(DWID - 1):0])
    ,.a_rid(split12_merge12_rid[(IDWID - 1):0])
    ,.a_rlast(split12_merge12_rlast)
    ,.a_rready(split12_merge12_rready)
    ,.a_rresp(split12_merge12_rresp[1:0])
    ,.a_rvalid(split12_merge12_rvalid)
    ,.a_wdata(split12_merge12_wdata[(DWID - 1):0])
    ,.a_wlast(split12_merge12_wlast)
    ,.a_wready(split12_merge12_wready)
    ,.a_wstrb(split12_merge12_wstrb[(WSTRB - 1):0])
    ,.a_wvalid(split12_merge12_wvalid)

    ,.b_araddr(split13_merge12_araddr[31:0])
    ,.b_arburst(split13_merge12_arburst[1:0])
    ,.b_arextras(split13_merge12_arextras[(EXTRAS - 1):0])
    ,.b_arid(split13_merge12_arid[(IDWID - 1):0])
    ,.b_arlen(split13_merge12_arlen[7:0])
    ,.b_arready(split13_merge12_arready)
    ,.b_arvalid(split13_merge12_arvalid)
    ,.b_awaddr(split13_merge12_awaddr[31:0])
    ,.b_awburst(split13_merge12_awburst[1:0])
    ,.b_awextras(split13_merge12_awextras[(EXTRAS - 1):0])
    ,.b_awid(split13_merge12_awid[(IDWID - 1):0])
    ,.b_awlen(split13_merge12_awlen[7:0])
    ,.b_awready(split13_merge12_awready)
    ,.b_awvalid(split13_merge12_awvalid)
    ,.b_bid(split13_merge12_bid[(IDWID - 1):0])
    ,.b_bready(split13_merge12_bready)
    ,.b_bresp(split13_merge12_bresp[1:0])
    ,.b_bvalid(split13_merge12_bvalid)
    ,.b_rdata(split13_merge12_rdata[(DWID - 1):0])
    ,.b_rid(split13_merge12_rid[(IDWID - 1):0])
    ,.b_rlast(split13_merge12_rlast)
    ,.b_rready(split13_merge12_rready)
    ,.b_rresp(split13_merge12_rresp[1:0])
    ,.b_rvalid(split13_merge12_rvalid)
    ,.b_wdata(split13_merge12_wdata[(DWID - 1):0])
    ,.b_wlast(split13_merge12_wlast)
    ,.b_wready(split13_merge12_wready)
    ,.b_wstrb(split13_merge12_wstrb[(WSTRB - 1):0])
    ,.b_wvalid(split13_merge12_wvalid)

    ,.c_araddr(split14_merge12_araddr[31:0])
    ,.c_arburst(split14_merge12_arburst[1:0])
    ,.c_arextras(split14_merge12_arextras[(EXTRAS - 1):0])
    ,.c_arid(split14_merge12_arid[(IDWID - 1):0])
    ,.c_arlen(split14_merge12_arlen[7:0])
    ,.c_arready(split14_merge12_arready)
    ,.c_arvalid(split14_merge12_arvalid)
    ,.c_awaddr(split14_merge12_awaddr[31:0])
    ,.c_awburst(split14_merge12_awburst[1:0])
    ,.c_awextras(split14_merge12_awextras[(EXTRAS - 1):0])
    ,.c_awid(split14_merge12_awid[(IDWID - 1):0])
    ,.c_awlen(split14_merge12_awlen[7:0])
    ,.c_awready(split14_merge12_awready)
    ,.c_awvalid(split14_merge12_awvalid)
    ,.c_bid(split14_merge12_bid[(IDWID - 1):0])
    ,.c_bready(split14_merge12_bready)
    ,.c_bresp(split14_merge12_bresp[1:0])
    ,.c_bvalid(split14_merge12_bvalid)
    ,.c_rdata(split14_merge12_rdata[(DWID - 1):0])
    ,.c_rid(split14_merge12_rid[(IDWID - 1):0])
    ,.c_rlast(split14_merge12_rlast)
    ,.c_rready(split14_merge12_rready)
    ,.c_rresp(split14_merge12_rresp[1:0])
    ,.c_rvalid(split14_merge12_rvalid)
    ,.c_wdata(split14_merge12_wdata[(DWID - 1):0])
    ,.c_wlast(split14_merge12_wlast)
    ,.c_wready(split14_merge12_wready)
    ,.c_wstrb(split14_merge12_wstrb[(WSTRB - 1):0])
    ,.c_wvalid(split14_merge12_wvalid)

    ,.d_araddr(split15_merge12_araddr[31:0])
    ,.d_arburst(split15_merge12_arburst[1:0])
    ,.d_arextras(split15_merge12_arextras[(EXTRAS - 1):0])
    ,.d_arid(split15_merge12_arid[(IDWID - 1):0])
    ,.d_arlen(split15_merge12_arlen[7:0])
    ,.d_arready(split15_merge12_arready)
    ,.d_arvalid(split15_merge12_arvalid)
    ,.d_awaddr(split15_merge12_awaddr[31:0])
    ,.d_awburst(split15_merge12_awburst[1:0])
    ,.d_awextras(split15_merge12_awextras[(EXTRAS - 1):0])
    ,.d_awid(split15_merge12_awid[(IDWID - 1):0])
    ,.d_awlen(split15_merge12_awlen[7:0])
    ,.d_awready(split15_merge12_awready)
    ,.d_awvalid(split15_merge12_awvalid)
    ,.d_bid(split15_merge12_bid[(IDWID - 1):0])
    ,.d_bready(split15_merge12_bready)
    ,.d_bresp(split15_merge12_bresp[1:0])
    ,.d_bvalid(split15_merge12_bvalid)
    ,.d_rdata(split15_merge12_rdata[(DWID - 1):0])
    ,.d_rid(split15_merge12_rid[(IDWID - 1):0])
    ,.d_rlast(split15_merge12_rlast)
    ,.d_rready(split15_merge12_rready)
    ,.d_rresp(split15_merge12_rresp[1:0])
    ,.d_rvalid(split15_merge12_rvalid)
    ,.d_wdata(split15_merge12_wdata[(DWID - 1):0])
    ,.d_wlast(split15_merge12_wlast)
    ,.d_wready(split15_merge12_wready)
    ,.d_wstrb(split15_merge12_wstrb[(WSTRB - 1):0])
    ,.d_wvalid(split15_merge12_wvalid)
);


wire [IDWID-1:0] merge13_split113_arid ;
wire [31:0] merge13_split113_araddr ;
wire [7:0] merge13_split113_arlen ;
wire [EXTRAS-1:0] merge13_split113_arextras ;
wire [1:0] merge13_split113_arburst ;
wire merge13_split113_arvalid ;
wire merge13_split113_arready ;
wire [IDWID-1:0] merge13_split113_rid ;
wire [DWID-1:0] merge13_split113_rdata ;
wire [1:0] merge13_split113_rresp ;
wire merge13_split113_rlast ;
wire merge13_split113_rvalid ;
wire merge13_split113_rready ;

wire [IDWID-1:0] merge13_split113_awid ;
wire [31:0] merge13_split113_awaddr ;
wire [7:0] merge13_split113_awlen ;
wire [EXTRAS-1:0] merge13_split113_awextras ;
wire [1:0] merge13_split113_awburst ;
wire merge13_split113_awvalid ;
wire merge13_split113_awready ;
wire [DWID-1:0] merge13_split113_wdata ;
wire [WSTRB-1:0] merge13_split113_wstrb ;
wire merge13_split113_wlast ;
wire merge13_split113_wvalid ;
wire merge13_split113_wready ;
wire [IDWID-1:0] merge13_split113_bid ;
wire [1:0] merge13_split113_bresp ;
wire merge13_split113_bvalid ;
wire merge13_split113_bready ;


wire [IDWID-1:0] split13_merge13_arid ;
wire [31:0] split13_merge13_araddr ;
wire [7:0] split13_merge13_arlen ;
wire [EXTRAS-1:0] split13_merge13_arextras ;
wire [1:0] split13_merge13_arburst ;
wire split13_merge13_arvalid ;
wire split13_merge13_arready ;
wire [IDWID-1:0] split13_merge13_rid ;
wire [DWID-1:0] split13_merge13_rdata ;
wire [1:0] split13_merge13_rresp ;
wire split13_merge13_rlast ;
wire split13_merge13_rvalid ;
wire split13_merge13_rready ;

wire [IDWID-1:0] split13_merge13_awid ;
wire [31:0] split13_merge13_awaddr ;
wire [7:0] split13_merge13_awlen ;
wire [EXTRAS-1:0] split13_merge13_awextras ;
wire [1:0] split13_merge13_awburst ;
wire split13_merge13_awvalid ;
wire split13_merge13_awready ;
wire [DWID-1:0] split13_merge13_wdata ;
wire [WSTRB-1:0] split13_merge13_wstrb ;
wire split13_merge13_wlast ;
wire split13_merge13_wvalid ;
wire split13_merge13_wready ;
wire [IDWID-1:0] split13_merge13_bid ;
wire [1:0] split13_merge13_bresp ;
wire split13_merge13_bvalid ;
wire split13_merge13_bready ;


wire [IDWID-1:0] split14_merge13_arid ;
wire [31:0] split14_merge13_araddr ;
wire [7:0] split14_merge13_arlen ;
wire [EXTRAS-1:0] split14_merge13_arextras ;
wire [1:0] split14_merge13_arburst ;
wire split14_merge13_arvalid ;
wire split14_merge13_arready ;
wire [IDWID-1:0] split14_merge13_rid ;
wire [DWID-1:0] split14_merge13_rdata ;
wire [1:0] split14_merge13_rresp ;
wire split14_merge13_rlast ;
wire split14_merge13_rvalid ;
wire split14_merge13_rready ;

wire [IDWID-1:0] split14_merge13_awid ;
wire [31:0] split14_merge13_awaddr ;
wire [7:0] split14_merge13_awlen ;
wire [EXTRAS-1:0] split14_merge13_awextras ;
wire [1:0] split14_merge13_awburst ;
wire split14_merge13_awvalid ;
wire split14_merge13_awready ;
wire [DWID-1:0] split14_merge13_wdata ;
wire [WSTRB-1:0] split14_merge13_wstrb ;
wire split14_merge13_wlast ;
wire split14_merge13_wvalid ;
wire split14_merge13_wready ;
wire [IDWID-1:0] split14_merge13_bid ;
wire [1:0] split14_merge13_bresp ;
wire split14_merge13_bvalid ;
wire split14_merge13_bready ;


wire [IDWID-1:0] split15_merge13_arid ;
wire [31:0] split15_merge13_araddr ;
wire [7:0] split15_merge13_arlen ;
wire [EXTRAS-1:0] split15_merge13_arextras ;
wire [1:0] split15_merge13_arburst ;
wire split15_merge13_arvalid ;
wire split15_merge13_arready ;
wire [IDWID-1:0] split15_merge13_rid ;
wire [DWID-1:0] split15_merge13_rdata ;
wire [1:0] split15_merge13_rresp ;
wire split15_merge13_rlast ;
wire split15_merge13_rvalid ;
wire split15_merge13_rready ;

wire [IDWID-1:0] split15_merge13_awid ;
wire [31:0] split15_merge13_awaddr ;
wire [7:0] split15_merge13_awlen ;
wire [EXTRAS-1:0] split15_merge13_awextras ;
wire [1:0] split15_merge13_awburst ;
wire split15_merge13_awvalid ;
wire split15_merge13_awready ;
wire [DWID-1:0] split15_merge13_wdata ;
wire [WSTRB-1:0] split15_merge13_wstrb ;
wire split15_merge13_wlast ;
wire split15_merge13_wvalid ;
wire split15_merge13_wready ;
wire [IDWID-1:0] split15_merge13_bid ;
wire [1:0] split15_merge13_bresp ;
wire split15_merge13_bvalid ;
wire split15_merge13_bready ;


axi_4_merger merge13 (
     .clk(clk),.rst_n(rst_n)
    ,.araddr(merge13_split113_araddr[31:0])
    ,.arburst(merge13_split113_arburst[1:0])
    ,.arextras(merge13_split113_arextras[(EXTRAS - 1):0])
    ,.arid(merge13_split113_arid[(IDWID - 1):0])
    ,.arlen(merge13_split113_arlen[7:0])
    ,.arready(merge13_split113_arready)
    ,.arvalid(merge13_split113_arvalid)
    ,.awaddr(merge13_split113_awaddr[31:0])
    ,.awburst(merge13_split113_awburst[1:0])
    ,.awextras(merge13_split113_awextras[(EXTRAS - 1):0])
    ,.awid(merge13_split113_awid[3:0])
    ,.awlen(merge13_split113_awlen[7:0])
    ,.awready(merge13_split113_awready)
    ,.awvalid(merge13_split113_awvalid)
    ,.bid(merge13_split113_bid[(IDWID - 1):0])
    ,.bready(merge13_split113_bready)
    ,.bresp(merge13_split113_bresp[1:0])
    ,.bvalid(merge13_split113_bvalid)
    ,.rid(merge13_split113_rid[(IDWID - 1):0])
    ,.rlast(merge13_split113_rlast)
    ,.rready(merge13_split113_rready)
    ,.rresp(merge13_split113_rresp[1:0])
    ,.rvalid(merge13_split113_rvalid)
    ,.rdata(merge13_split113_rdata[(DWID - 1):0])
    ,.wdata(merge13_split113_wdata[(DWID - 1):0])
    ,.wlast(merge13_split113_wlast)
    ,.wready(merge13_split113_wready)
    ,.wstrb(merge13_split113_wstrb[(WSTRB - 1):0])
    ,.wvalid(merge13_split113_wvalid)


    ,.a_araddr(split12_merge13_araddr[31:0])
    ,.a_arburst(split12_merge13_arburst[1:0])
    ,.a_arextras(split12_merge13_arextras[(EXTRAS - 1):0])
    ,.a_arid(split12_merge13_arid[(IDWID - 1):0])
    ,.a_arlen(split12_merge13_arlen[7:0])
    ,.a_arready(split12_merge13_arready)
    ,.a_arvalid(split12_merge13_arvalid)
    ,.a_awaddr(split12_merge13_awaddr[31:0])
    ,.a_awburst(split12_merge13_awburst[1:0])
    ,.a_awextras(split12_merge13_awextras[(EXTRAS - 1):0])
    ,.a_awid(split12_merge13_awid[(IDWID - 1):0])
    ,.a_awlen(split12_merge13_awlen[7:0])
    ,.a_awready(split12_merge13_awready)
    ,.a_awvalid(split12_merge13_awvalid)
    ,.a_bid(split12_merge13_bid[(IDWID - 1):0])
    ,.a_bready(split12_merge13_bready)
    ,.a_bresp(split12_merge13_bresp[1:0])
    ,.a_bvalid(split12_merge13_bvalid)
    ,.a_rdata(split12_merge13_rdata[(DWID - 1):0])
    ,.a_rid(split12_merge13_rid[(IDWID - 1):0])
    ,.a_rlast(split12_merge13_rlast)
    ,.a_rready(split12_merge13_rready)
    ,.a_rresp(split12_merge13_rresp[1:0])
    ,.a_rvalid(split12_merge13_rvalid)
    ,.a_wdata(split12_merge13_wdata[(DWID - 1):0])
    ,.a_wlast(split12_merge13_wlast)
    ,.a_wready(split12_merge13_wready)
    ,.a_wstrb(split12_merge13_wstrb[(WSTRB - 1):0])
    ,.a_wvalid(split12_merge13_wvalid)

    ,.b_araddr(split13_merge13_araddr[31:0])
    ,.b_arburst(split13_merge13_arburst[1:0])
    ,.b_arextras(split13_merge13_arextras[(EXTRAS - 1):0])
    ,.b_arid(split13_merge13_arid[(IDWID - 1):0])
    ,.b_arlen(split13_merge13_arlen[7:0])
    ,.b_arready(split13_merge13_arready)
    ,.b_arvalid(split13_merge13_arvalid)
    ,.b_awaddr(split13_merge13_awaddr[31:0])
    ,.b_awburst(split13_merge13_awburst[1:0])
    ,.b_awextras(split13_merge13_awextras[(EXTRAS - 1):0])
    ,.b_awid(split13_merge13_awid[(IDWID - 1):0])
    ,.b_awlen(split13_merge13_awlen[7:0])
    ,.b_awready(split13_merge13_awready)
    ,.b_awvalid(split13_merge13_awvalid)
    ,.b_bid(split13_merge13_bid[(IDWID - 1):0])
    ,.b_bready(split13_merge13_bready)
    ,.b_bresp(split13_merge13_bresp[1:0])
    ,.b_bvalid(split13_merge13_bvalid)
    ,.b_rdata(split13_merge13_rdata[(DWID - 1):0])
    ,.b_rid(split13_merge13_rid[(IDWID - 1):0])
    ,.b_rlast(split13_merge13_rlast)
    ,.b_rready(split13_merge13_rready)
    ,.b_rresp(split13_merge13_rresp[1:0])
    ,.b_rvalid(split13_merge13_rvalid)
    ,.b_wdata(split13_merge13_wdata[(DWID - 1):0])
    ,.b_wlast(split13_merge13_wlast)
    ,.b_wready(split13_merge13_wready)
    ,.b_wstrb(split13_merge13_wstrb[(WSTRB - 1):0])
    ,.b_wvalid(split13_merge13_wvalid)

    ,.c_araddr(split14_merge13_araddr[31:0])
    ,.c_arburst(split14_merge13_arburst[1:0])
    ,.c_arextras(split14_merge13_arextras[(EXTRAS - 1):0])
    ,.c_arid(split14_merge13_arid[(IDWID - 1):0])
    ,.c_arlen(split14_merge13_arlen[7:0])
    ,.c_arready(split14_merge13_arready)
    ,.c_arvalid(split14_merge13_arvalid)
    ,.c_awaddr(split14_merge13_awaddr[31:0])
    ,.c_awburst(split14_merge13_awburst[1:0])
    ,.c_awextras(split14_merge13_awextras[(EXTRAS - 1):0])
    ,.c_awid(split14_merge13_awid[(IDWID - 1):0])
    ,.c_awlen(split14_merge13_awlen[7:0])
    ,.c_awready(split14_merge13_awready)
    ,.c_awvalid(split14_merge13_awvalid)
    ,.c_bid(split14_merge13_bid[(IDWID - 1):0])
    ,.c_bready(split14_merge13_bready)
    ,.c_bresp(split14_merge13_bresp[1:0])
    ,.c_bvalid(split14_merge13_bvalid)
    ,.c_rdata(split14_merge13_rdata[(DWID - 1):0])
    ,.c_rid(split14_merge13_rid[(IDWID - 1):0])
    ,.c_rlast(split14_merge13_rlast)
    ,.c_rready(split14_merge13_rready)
    ,.c_rresp(split14_merge13_rresp[1:0])
    ,.c_rvalid(split14_merge13_rvalid)
    ,.c_wdata(split14_merge13_wdata[(DWID - 1):0])
    ,.c_wlast(split14_merge13_wlast)
    ,.c_wready(split14_merge13_wready)
    ,.c_wstrb(split14_merge13_wstrb[(WSTRB - 1):0])
    ,.c_wvalid(split14_merge13_wvalid)

    ,.d_araddr(split15_merge13_araddr[31:0])
    ,.d_arburst(split15_merge13_arburst[1:0])
    ,.d_arextras(split15_merge13_arextras[(EXTRAS - 1):0])
    ,.d_arid(split15_merge13_arid[(IDWID - 1):0])
    ,.d_arlen(split15_merge13_arlen[7:0])
    ,.d_arready(split15_merge13_arready)
    ,.d_arvalid(split15_merge13_arvalid)
    ,.d_awaddr(split15_merge13_awaddr[31:0])
    ,.d_awburst(split15_merge13_awburst[1:0])
    ,.d_awextras(split15_merge13_awextras[(EXTRAS - 1):0])
    ,.d_awid(split15_merge13_awid[(IDWID - 1):0])
    ,.d_awlen(split15_merge13_awlen[7:0])
    ,.d_awready(split15_merge13_awready)
    ,.d_awvalid(split15_merge13_awvalid)
    ,.d_bid(split15_merge13_bid[(IDWID - 1):0])
    ,.d_bready(split15_merge13_bready)
    ,.d_bresp(split15_merge13_bresp[1:0])
    ,.d_bvalid(split15_merge13_bvalid)
    ,.d_rdata(split15_merge13_rdata[(DWID - 1):0])
    ,.d_rid(split15_merge13_rid[(IDWID - 1):0])
    ,.d_rlast(split15_merge13_rlast)
    ,.d_rready(split15_merge13_rready)
    ,.d_rresp(split15_merge13_rresp[1:0])
    ,.d_rvalid(split15_merge13_rvalid)
    ,.d_wdata(split15_merge13_wdata[(DWID - 1):0])
    ,.d_wlast(split15_merge13_wlast)
    ,.d_wready(split15_merge13_wready)
    ,.d_wstrb(split15_merge13_wstrb[(WSTRB - 1):0])
    ,.d_wvalid(split15_merge13_wvalid)
);


wire [IDWID-1:0] merge14_split114_arid ;
wire [31:0] merge14_split114_araddr ;
wire [7:0] merge14_split114_arlen ;
wire [EXTRAS-1:0] merge14_split114_arextras ;
wire [1:0] merge14_split114_arburst ;
wire merge14_split114_arvalid ;
wire merge14_split114_arready ;
wire [IDWID-1:0] merge14_split114_rid ;
wire [DWID-1:0] merge14_split114_rdata ;
wire [1:0] merge14_split114_rresp ;
wire merge14_split114_rlast ;
wire merge14_split114_rvalid ;
wire merge14_split114_rready ;

wire [IDWID-1:0] merge14_split114_awid ;
wire [31:0] merge14_split114_awaddr ;
wire [7:0] merge14_split114_awlen ;
wire [EXTRAS-1:0] merge14_split114_awextras ;
wire [1:0] merge14_split114_awburst ;
wire merge14_split114_awvalid ;
wire merge14_split114_awready ;
wire [DWID-1:0] merge14_split114_wdata ;
wire [WSTRB-1:0] merge14_split114_wstrb ;
wire merge14_split114_wlast ;
wire merge14_split114_wvalid ;
wire merge14_split114_wready ;
wire [IDWID-1:0] merge14_split114_bid ;
wire [1:0] merge14_split114_bresp ;
wire merge14_split114_bvalid ;
wire merge14_split114_bready ;


wire [IDWID-1:0] split13_merge14_arid ;
wire [31:0] split13_merge14_araddr ;
wire [7:0] split13_merge14_arlen ;
wire [EXTRAS-1:0] split13_merge14_arextras ;
wire [1:0] split13_merge14_arburst ;
wire split13_merge14_arvalid ;
wire split13_merge14_arready ;
wire [IDWID-1:0] split13_merge14_rid ;
wire [DWID-1:0] split13_merge14_rdata ;
wire [1:0] split13_merge14_rresp ;
wire split13_merge14_rlast ;
wire split13_merge14_rvalid ;
wire split13_merge14_rready ;

wire [IDWID-1:0] split13_merge14_awid ;
wire [31:0] split13_merge14_awaddr ;
wire [7:0] split13_merge14_awlen ;
wire [EXTRAS-1:0] split13_merge14_awextras ;
wire [1:0] split13_merge14_awburst ;
wire split13_merge14_awvalid ;
wire split13_merge14_awready ;
wire [DWID-1:0] split13_merge14_wdata ;
wire [WSTRB-1:0] split13_merge14_wstrb ;
wire split13_merge14_wlast ;
wire split13_merge14_wvalid ;
wire split13_merge14_wready ;
wire [IDWID-1:0] split13_merge14_bid ;
wire [1:0] split13_merge14_bresp ;
wire split13_merge14_bvalid ;
wire split13_merge14_bready ;


wire [IDWID-1:0] split14_merge14_arid ;
wire [31:0] split14_merge14_araddr ;
wire [7:0] split14_merge14_arlen ;
wire [EXTRAS-1:0] split14_merge14_arextras ;
wire [1:0] split14_merge14_arburst ;
wire split14_merge14_arvalid ;
wire split14_merge14_arready ;
wire [IDWID-1:0] split14_merge14_rid ;
wire [DWID-1:0] split14_merge14_rdata ;
wire [1:0] split14_merge14_rresp ;
wire split14_merge14_rlast ;
wire split14_merge14_rvalid ;
wire split14_merge14_rready ;

wire [IDWID-1:0] split14_merge14_awid ;
wire [31:0] split14_merge14_awaddr ;
wire [7:0] split14_merge14_awlen ;
wire [EXTRAS-1:0] split14_merge14_awextras ;
wire [1:0] split14_merge14_awburst ;
wire split14_merge14_awvalid ;
wire split14_merge14_awready ;
wire [DWID-1:0] split14_merge14_wdata ;
wire [WSTRB-1:0] split14_merge14_wstrb ;
wire split14_merge14_wlast ;
wire split14_merge14_wvalid ;
wire split14_merge14_wready ;
wire [IDWID-1:0] split14_merge14_bid ;
wire [1:0] split14_merge14_bresp ;
wire split14_merge14_bvalid ;
wire split14_merge14_bready ;


wire [IDWID-1:0] split15_merge14_arid ;
wire [31:0] split15_merge14_araddr ;
wire [7:0] split15_merge14_arlen ;
wire [EXTRAS-1:0] split15_merge14_arextras ;
wire [1:0] split15_merge14_arburst ;
wire split15_merge14_arvalid ;
wire split15_merge14_arready ;
wire [IDWID-1:0] split15_merge14_rid ;
wire [DWID-1:0] split15_merge14_rdata ;
wire [1:0] split15_merge14_rresp ;
wire split15_merge14_rlast ;
wire split15_merge14_rvalid ;
wire split15_merge14_rready ;

wire [IDWID-1:0] split15_merge14_awid ;
wire [31:0] split15_merge14_awaddr ;
wire [7:0] split15_merge14_awlen ;
wire [EXTRAS-1:0] split15_merge14_awextras ;
wire [1:0] split15_merge14_awburst ;
wire split15_merge14_awvalid ;
wire split15_merge14_awready ;
wire [DWID-1:0] split15_merge14_wdata ;
wire [WSTRB-1:0] split15_merge14_wstrb ;
wire split15_merge14_wlast ;
wire split15_merge14_wvalid ;
wire split15_merge14_wready ;
wire [IDWID-1:0] split15_merge14_bid ;
wire [1:0] split15_merge14_bresp ;
wire split15_merge14_bvalid ;
wire split15_merge14_bready ;


axi_4_merger merge14 (
     .clk(clk),.rst_n(rst_n)
    ,.araddr(merge14_split114_araddr[31:0])
    ,.arburst(merge14_split114_arburst[1:0])
    ,.arextras(merge14_split114_arextras[(EXTRAS - 1):0])
    ,.arid(merge14_split114_arid[(IDWID - 1):0])
    ,.arlen(merge14_split114_arlen[7:0])
    ,.arready(merge14_split114_arready)
    ,.arvalid(merge14_split114_arvalid)
    ,.awaddr(merge14_split114_awaddr[31:0])
    ,.awburst(merge14_split114_awburst[1:0])
    ,.awextras(merge14_split114_awextras[(EXTRAS - 1):0])
    ,.awid(merge14_split114_awid[3:0])
    ,.awlen(merge14_split114_awlen[7:0])
    ,.awready(merge14_split114_awready)
    ,.awvalid(merge14_split114_awvalid)
    ,.bid(merge14_split114_bid[(IDWID - 1):0])
    ,.bready(merge14_split114_bready)
    ,.bresp(merge14_split114_bresp[1:0])
    ,.bvalid(merge14_split114_bvalid)
    ,.rid(merge14_split114_rid[(IDWID - 1):0])
    ,.rlast(merge14_split114_rlast)
    ,.rready(merge14_split114_rready)
    ,.rresp(merge14_split114_rresp[1:0])
    ,.rvalid(merge14_split114_rvalid)
    ,.rdata(merge14_split114_rdata[(DWID - 1):0])
    ,.wdata(merge14_split114_wdata[(DWID - 1):0])
    ,.wlast(merge14_split114_wlast)
    ,.wready(merge14_split114_wready)
    ,.wstrb(merge14_split114_wstrb[(WSTRB - 1):0])
    ,.wvalid(merge14_split114_wvalid)


    ,.a_araddr(split12_merge14_araddr[31:0])
    ,.a_arburst(split12_merge14_arburst[1:0])
    ,.a_arextras(split12_merge14_arextras[(EXTRAS - 1):0])
    ,.a_arid(split12_merge14_arid[(IDWID - 1):0])
    ,.a_arlen(split12_merge14_arlen[7:0])
    ,.a_arready(split12_merge14_arready)
    ,.a_arvalid(split12_merge14_arvalid)
    ,.a_awaddr(split12_merge14_awaddr[31:0])
    ,.a_awburst(split12_merge14_awburst[1:0])
    ,.a_awextras(split12_merge14_awextras[(EXTRAS - 1):0])
    ,.a_awid(split12_merge14_awid[(IDWID - 1):0])
    ,.a_awlen(split12_merge14_awlen[7:0])
    ,.a_awready(split12_merge14_awready)
    ,.a_awvalid(split12_merge14_awvalid)
    ,.a_bid(split12_merge14_bid[(IDWID - 1):0])
    ,.a_bready(split12_merge14_bready)
    ,.a_bresp(split12_merge14_bresp[1:0])
    ,.a_bvalid(split12_merge14_bvalid)
    ,.a_rdata(split12_merge14_rdata[(DWID - 1):0])
    ,.a_rid(split12_merge14_rid[(IDWID - 1):0])
    ,.a_rlast(split12_merge14_rlast)
    ,.a_rready(split12_merge14_rready)
    ,.a_rresp(split12_merge14_rresp[1:0])
    ,.a_rvalid(split12_merge14_rvalid)
    ,.a_wdata(split12_merge14_wdata[(DWID - 1):0])
    ,.a_wlast(split12_merge14_wlast)
    ,.a_wready(split12_merge14_wready)
    ,.a_wstrb(split12_merge14_wstrb[(WSTRB - 1):0])
    ,.a_wvalid(split12_merge14_wvalid)

    ,.b_araddr(split13_merge14_araddr[31:0])
    ,.b_arburst(split13_merge14_arburst[1:0])
    ,.b_arextras(split13_merge14_arextras[(EXTRAS - 1):0])
    ,.b_arid(split13_merge14_arid[(IDWID - 1):0])
    ,.b_arlen(split13_merge14_arlen[7:0])
    ,.b_arready(split13_merge14_arready)
    ,.b_arvalid(split13_merge14_arvalid)
    ,.b_awaddr(split13_merge14_awaddr[31:0])
    ,.b_awburst(split13_merge14_awburst[1:0])
    ,.b_awextras(split13_merge14_awextras[(EXTRAS - 1):0])
    ,.b_awid(split13_merge14_awid[(IDWID - 1):0])
    ,.b_awlen(split13_merge14_awlen[7:0])
    ,.b_awready(split13_merge14_awready)
    ,.b_awvalid(split13_merge14_awvalid)
    ,.b_bid(split13_merge14_bid[(IDWID - 1):0])
    ,.b_bready(split13_merge14_bready)
    ,.b_bresp(split13_merge14_bresp[1:0])
    ,.b_bvalid(split13_merge14_bvalid)
    ,.b_rdata(split13_merge14_rdata[(DWID - 1):0])
    ,.b_rid(split13_merge14_rid[(IDWID - 1):0])
    ,.b_rlast(split13_merge14_rlast)
    ,.b_rready(split13_merge14_rready)
    ,.b_rresp(split13_merge14_rresp[1:0])
    ,.b_rvalid(split13_merge14_rvalid)
    ,.b_wdata(split13_merge14_wdata[(DWID - 1):0])
    ,.b_wlast(split13_merge14_wlast)
    ,.b_wready(split13_merge14_wready)
    ,.b_wstrb(split13_merge14_wstrb[(WSTRB - 1):0])
    ,.b_wvalid(split13_merge14_wvalid)

    ,.c_araddr(split14_merge14_araddr[31:0])
    ,.c_arburst(split14_merge14_arburst[1:0])
    ,.c_arextras(split14_merge14_arextras[(EXTRAS - 1):0])
    ,.c_arid(split14_merge14_arid[(IDWID - 1):0])
    ,.c_arlen(split14_merge14_arlen[7:0])
    ,.c_arready(split14_merge14_arready)
    ,.c_arvalid(split14_merge14_arvalid)
    ,.c_awaddr(split14_merge14_awaddr[31:0])
    ,.c_awburst(split14_merge14_awburst[1:0])
    ,.c_awextras(split14_merge14_awextras[(EXTRAS - 1):0])
    ,.c_awid(split14_merge14_awid[(IDWID - 1):0])
    ,.c_awlen(split14_merge14_awlen[7:0])
    ,.c_awready(split14_merge14_awready)
    ,.c_awvalid(split14_merge14_awvalid)
    ,.c_bid(split14_merge14_bid[(IDWID - 1):0])
    ,.c_bready(split14_merge14_bready)
    ,.c_bresp(split14_merge14_bresp[1:0])
    ,.c_bvalid(split14_merge14_bvalid)
    ,.c_rdata(split14_merge14_rdata[(DWID - 1):0])
    ,.c_rid(split14_merge14_rid[(IDWID - 1):0])
    ,.c_rlast(split14_merge14_rlast)
    ,.c_rready(split14_merge14_rready)
    ,.c_rresp(split14_merge14_rresp[1:0])
    ,.c_rvalid(split14_merge14_rvalid)
    ,.c_wdata(split14_merge14_wdata[(DWID - 1):0])
    ,.c_wlast(split14_merge14_wlast)
    ,.c_wready(split14_merge14_wready)
    ,.c_wstrb(split14_merge14_wstrb[(WSTRB - 1):0])
    ,.c_wvalid(split14_merge14_wvalid)

    ,.d_araddr(split15_merge14_araddr[31:0])
    ,.d_arburst(split15_merge14_arburst[1:0])
    ,.d_arextras(split15_merge14_arextras[(EXTRAS - 1):0])
    ,.d_arid(split15_merge14_arid[(IDWID - 1):0])
    ,.d_arlen(split15_merge14_arlen[7:0])
    ,.d_arready(split15_merge14_arready)
    ,.d_arvalid(split15_merge14_arvalid)
    ,.d_awaddr(split15_merge14_awaddr[31:0])
    ,.d_awburst(split15_merge14_awburst[1:0])
    ,.d_awextras(split15_merge14_awextras[(EXTRAS - 1):0])
    ,.d_awid(split15_merge14_awid[(IDWID - 1):0])
    ,.d_awlen(split15_merge14_awlen[7:0])
    ,.d_awready(split15_merge14_awready)
    ,.d_awvalid(split15_merge14_awvalid)
    ,.d_bid(split15_merge14_bid[(IDWID - 1):0])
    ,.d_bready(split15_merge14_bready)
    ,.d_bresp(split15_merge14_bresp[1:0])
    ,.d_bvalid(split15_merge14_bvalid)
    ,.d_rdata(split15_merge14_rdata[(DWID - 1):0])
    ,.d_rid(split15_merge14_rid[(IDWID - 1):0])
    ,.d_rlast(split15_merge14_rlast)
    ,.d_rready(split15_merge14_rready)
    ,.d_rresp(split15_merge14_rresp[1:0])
    ,.d_rvalid(split15_merge14_rvalid)
    ,.d_wdata(split15_merge14_wdata[(DWID - 1):0])
    ,.d_wlast(split15_merge14_wlast)
    ,.d_wready(split15_merge14_wready)
    ,.d_wstrb(split15_merge14_wstrb[(WSTRB - 1):0])
    ,.d_wvalid(split15_merge14_wvalid)
);


wire [IDWID-1:0] merge15_split115_arid ;
wire [31:0] merge15_split115_araddr ;
wire [7:0] merge15_split115_arlen ;
wire [EXTRAS-1:0] merge15_split115_arextras ;
wire [1:0] merge15_split115_arburst ;
wire merge15_split115_arvalid ;
wire merge15_split115_arready ;
wire [IDWID-1:0] merge15_split115_rid ;
wire [DWID-1:0] merge15_split115_rdata ;
wire [1:0] merge15_split115_rresp ;
wire merge15_split115_rlast ;
wire merge15_split115_rvalid ;
wire merge15_split115_rready ;

wire [IDWID-1:0] merge15_split115_awid ;
wire [31:0] merge15_split115_awaddr ;
wire [7:0] merge15_split115_awlen ;
wire [EXTRAS-1:0] merge15_split115_awextras ;
wire [1:0] merge15_split115_awburst ;
wire merge15_split115_awvalid ;
wire merge15_split115_awready ;
wire [DWID-1:0] merge15_split115_wdata ;
wire [WSTRB-1:0] merge15_split115_wstrb ;
wire merge15_split115_wlast ;
wire merge15_split115_wvalid ;
wire merge15_split115_wready ;
wire [IDWID-1:0] merge15_split115_bid ;
wire [1:0] merge15_split115_bresp ;
wire merge15_split115_bvalid ;
wire merge15_split115_bready ;


wire [IDWID-1:0] split13_merge15_arid ;
wire [31:0] split13_merge15_araddr ;
wire [7:0] split13_merge15_arlen ;
wire [EXTRAS-1:0] split13_merge15_arextras ;
wire [1:0] split13_merge15_arburst ;
wire split13_merge15_arvalid ;
wire split13_merge15_arready ;
wire [IDWID-1:0] split13_merge15_rid ;
wire [DWID-1:0] split13_merge15_rdata ;
wire [1:0] split13_merge15_rresp ;
wire split13_merge15_rlast ;
wire split13_merge15_rvalid ;
wire split13_merge15_rready ;

wire [IDWID-1:0] split13_merge15_awid ;
wire [31:0] split13_merge15_awaddr ;
wire [7:0] split13_merge15_awlen ;
wire [EXTRAS-1:0] split13_merge15_awextras ;
wire [1:0] split13_merge15_awburst ;
wire split13_merge15_awvalid ;
wire split13_merge15_awready ;
wire [DWID-1:0] split13_merge15_wdata ;
wire [WSTRB-1:0] split13_merge15_wstrb ;
wire split13_merge15_wlast ;
wire split13_merge15_wvalid ;
wire split13_merge15_wready ;
wire [IDWID-1:0] split13_merge15_bid ;
wire [1:0] split13_merge15_bresp ;
wire split13_merge15_bvalid ;
wire split13_merge15_bready ;


wire [IDWID-1:0] split14_merge15_arid ;
wire [31:0] split14_merge15_araddr ;
wire [7:0] split14_merge15_arlen ;
wire [EXTRAS-1:0] split14_merge15_arextras ;
wire [1:0] split14_merge15_arburst ;
wire split14_merge15_arvalid ;
wire split14_merge15_arready ;
wire [IDWID-1:0] split14_merge15_rid ;
wire [DWID-1:0] split14_merge15_rdata ;
wire [1:0] split14_merge15_rresp ;
wire split14_merge15_rlast ;
wire split14_merge15_rvalid ;
wire split14_merge15_rready ;

wire [IDWID-1:0] split14_merge15_awid ;
wire [31:0] split14_merge15_awaddr ;
wire [7:0] split14_merge15_awlen ;
wire [EXTRAS-1:0] split14_merge15_awextras ;
wire [1:0] split14_merge15_awburst ;
wire split14_merge15_awvalid ;
wire split14_merge15_awready ;
wire [DWID-1:0] split14_merge15_wdata ;
wire [WSTRB-1:0] split14_merge15_wstrb ;
wire split14_merge15_wlast ;
wire split14_merge15_wvalid ;
wire split14_merge15_wready ;
wire [IDWID-1:0] split14_merge15_bid ;
wire [1:0] split14_merge15_bresp ;
wire split14_merge15_bvalid ;
wire split14_merge15_bready ;


wire [IDWID-1:0] split15_merge15_arid ;
wire [31:0] split15_merge15_araddr ;
wire [7:0] split15_merge15_arlen ;
wire [EXTRAS-1:0] split15_merge15_arextras ;
wire [1:0] split15_merge15_arburst ;
wire split15_merge15_arvalid ;
wire split15_merge15_arready ;
wire [IDWID-1:0] split15_merge15_rid ;
wire [DWID-1:0] split15_merge15_rdata ;
wire [1:0] split15_merge15_rresp ;
wire split15_merge15_rlast ;
wire split15_merge15_rvalid ;
wire split15_merge15_rready ;

wire [IDWID-1:0] split15_merge15_awid ;
wire [31:0] split15_merge15_awaddr ;
wire [7:0] split15_merge15_awlen ;
wire [EXTRAS-1:0] split15_merge15_awextras ;
wire [1:0] split15_merge15_awburst ;
wire split15_merge15_awvalid ;
wire split15_merge15_awready ;
wire [DWID-1:0] split15_merge15_wdata ;
wire [WSTRB-1:0] split15_merge15_wstrb ;
wire split15_merge15_wlast ;
wire split15_merge15_wvalid ;
wire split15_merge15_wready ;
wire [IDWID-1:0] split15_merge15_bid ;
wire [1:0] split15_merge15_bresp ;
wire split15_merge15_bvalid ;
wire split15_merge15_bready ;


axi_4_merger merge15 (
     .clk(clk),.rst_n(rst_n)
    ,.araddr(merge15_split115_araddr[31:0])
    ,.arburst(merge15_split115_arburst[1:0])
    ,.arextras(merge15_split115_arextras[(EXTRAS - 1):0])
    ,.arid(merge15_split115_arid[(IDWID - 1):0])
    ,.arlen(merge15_split115_arlen[7:0])
    ,.arready(merge15_split115_arready)
    ,.arvalid(merge15_split115_arvalid)
    ,.awaddr(merge15_split115_awaddr[31:0])
    ,.awburst(merge15_split115_awburst[1:0])
    ,.awextras(merge15_split115_awextras[(EXTRAS - 1):0])
    ,.awid(merge15_split115_awid[3:0])
    ,.awlen(merge15_split115_awlen[7:0])
    ,.awready(merge15_split115_awready)
    ,.awvalid(merge15_split115_awvalid)
    ,.bid(merge15_split115_bid[(IDWID - 1):0])
    ,.bready(merge15_split115_bready)
    ,.bresp(merge15_split115_bresp[1:0])
    ,.bvalid(merge15_split115_bvalid)
    ,.rid(merge15_split115_rid[(IDWID - 1):0])
    ,.rlast(merge15_split115_rlast)
    ,.rready(merge15_split115_rready)
    ,.rresp(merge15_split115_rresp[1:0])
    ,.rvalid(merge15_split115_rvalid)
    ,.rdata(merge15_split115_rdata[(DWID - 1):0])
    ,.wdata(merge15_split115_wdata[(DWID - 1):0])
    ,.wlast(merge15_split115_wlast)
    ,.wready(merge15_split115_wready)
    ,.wstrb(merge15_split115_wstrb[(WSTRB - 1):0])
    ,.wvalid(merge15_split115_wvalid)


    ,.a_araddr(split12_merge15_araddr[31:0])
    ,.a_arburst(split12_merge15_arburst[1:0])
    ,.a_arextras(split12_merge15_arextras[(EXTRAS - 1):0])
    ,.a_arid(split12_merge15_arid[(IDWID - 1):0])
    ,.a_arlen(split12_merge15_arlen[7:0])
    ,.a_arready(split12_merge15_arready)
    ,.a_arvalid(split12_merge15_arvalid)
    ,.a_awaddr(split12_merge15_awaddr[31:0])
    ,.a_awburst(split12_merge15_awburst[1:0])
    ,.a_awextras(split12_merge15_awextras[(EXTRAS - 1):0])
    ,.a_awid(split12_merge15_awid[(IDWID - 1):0])
    ,.a_awlen(split12_merge15_awlen[7:0])
    ,.a_awready(split12_merge15_awready)
    ,.a_awvalid(split12_merge15_awvalid)
    ,.a_bid(split12_merge15_bid[(IDWID - 1):0])
    ,.a_bready(split12_merge15_bready)
    ,.a_bresp(split12_merge15_bresp[1:0])
    ,.a_bvalid(split12_merge15_bvalid)
    ,.a_rdata(split12_merge15_rdata[(DWID - 1):0])
    ,.a_rid(split12_merge15_rid[(IDWID - 1):0])
    ,.a_rlast(split12_merge15_rlast)
    ,.a_rready(split12_merge15_rready)
    ,.a_rresp(split12_merge15_rresp[1:0])
    ,.a_rvalid(split12_merge15_rvalid)
    ,.a_wdata(split12_merge15_wdata[(DWID - 1):0])
    ,.a_wlast(split12_merge15_wlast)
    ,.a_wready(split12_merge15_wready)
    ,.a_wstrb(split12_merge15_wstrb[(WSTRB - 1):0])
    ,.a_wvalid(split12_merge15_wvalid)

    ,.b_araddr(split13_merge15_araddr[31:0])
    ,.b_arburst(split13_merge15_arburst[1:0])
    ,.b_arextras(split13_merge15_arextras[(EXTRAS - 1):0])
    ,.b_arid(split13_merge15_arid[(IDWID - 1):0])
    ,.b_arlen(split13_merge15_arlen[7:0])
    ,.b_arready(split13_merge15_arready)
    ,.b_arvalid(split13_merge15_arvalid)
    ,.b_awaddr(split13_merge15_awaddr[31:0])
    ,.b_awburst(split13_merge15_awburst[1:0])
    ,.b_awextras(split13_merge15_awextras[(EXTRAS - 1):0])
    ,.b_awid(split13_merge15_awid[(IDWID - 1):0])
    ,.b_awlen(split13_merge15_awlen[7:0])
    ,.b_awready(split13_merge15_awready)
    ,.b_awvalid(split13_merge15_awvalid)
    ,.b_bid(split13_merge15_bid[(IDWID - 1):0])
    ,.b_bready(split13_merge15_bready)
    ,.b_bresp(split13_merge15_bresp[1:0])
    ,.b_bvalid(split13_merge15_bvalid)
    ,.b_rdata(split13_merge15_rdata[(DWID - 1):0])
    ,.b_rid(split13_merge15_rid[(IDWID - 1):0])
    ,.b_rlast(split13_merge15_rlast)
    ,.b_rready(split13_merge15_rready)
    ,.b_rresp(split13_merge15_rresp[1:0])
    ,.b_rvalid(split13_merge15_rvalid)
    ,.b_wdata(split13_merge15_wdata[(DWID - 1):0])
    ,.b_wlast(split13_merge15_wlast)
    ,.b_wready(split13_merge15_wready)
    ,.b_wstrb(split13_merge15_wstrb[(WSTRB - 1):0])
    ,.b_wvalid(split13_merge15_wvalid)

    ,.c_araddr(split14_merge15_araddr[31:0])
    ,.c_arburst(split14_merge15_arburst[1:0])
    ,.c_arextras(split14_merge15_arextras[(EXTRAS - 1):0])
    ,.c_arid(split14_merge15_arid[(IDWID - 1):0])
    ,.c_arlen(split14_merge15_arlen[7:0])
    ,.c_arready(split14_merge15_arready)
    ,.c_arvalid(split14_merge15_arvalid)
    ,.c_awaddr(split14_merge15_awaddr[31:0])
    ,.c_awburst(split14_merge15_awburst[1:0])
    ,.c_awextras(split14_merge15_awextras[(EXTRAS - 1):0])
    ,.c_awid(split14_merge15_awid[(IDWID - 1):0])
    ,.c_awlen(split14_merge15_awlen[7:0])
    ,.c_awready(split14_merge15_awready)
    ,.c_awvalid(split14_merge15_awvalid)
    ,.c_bid(split14_merge15_bid[(IDWID - 1):0])
    ,.c_bready(split14_merge15_bready)
    ,.c_bresp(split14_merge15_bresp[1:0])
    ,.c_bvalid(split14_merge15_bvalid)
    ,.c_rdata(split14_merge15_rdata[(DWID - 1):0])
    ,.c_rid(split14_merge15_rid[(IDWID - 1):0])
    ,.c_rlast(split14_merge15_rlast)
    ,.c_rready(split14_merge15_rready)
    ,.c_rresp(split14_merge15_rresp[1:0])
    ,.c_rvalid(split14_merge15_rvalid)
    ,.c_wdata(split14_merge15_wdata[(DWID - 1):0])
    ,.c_wlast(split14_merge15_wlast)
    ,.c_wready(split14_merge15_wready)
    ,.c_wstrb(split14_merge15_wstrb[(WSTRB - 1):0])
    ,.c_wvalid(split14_merge15_wvalid)

    ,.d_araddr(split15_merge15_araddr[31:0])
    ,.d_arburst(split15_merge15_arburst[1:0])
    ,.d_arextras(split15_merge15_arextras[(EXTRAS - 1):0])
    ,.d_arid(split15_merge15_arid[(IDWID - 1):0])
    ,.d_arlen(split15_merge15_arlen[7:0])
    ,.d_arready(split15_merge15_arready)
    ,.d_arvalid(split15_merge15_arvalid)
    ,.d_awaddr(split15_merge15_awaddr[31:0])
    ,.d_awburst(split15_merge15_awburst[1:0])
    ,.d_awextras(split15_merge15_awextras[(EXTRAS - 1):0])
    ,.d_awid(split15_merge15_awid[(IDWID - 1):0])
    ,.d_awlen(split15_merge15_awlen[7:0])
    ,.d_awready(split15_merge15_awready)
    ,.d_awvalid(split15_merge15_awvalid)
    ,.d_bid(split15_merge15_bid[(IDWID - 1):0])
    ,.d_bready(split15_merge15_bready)
    ,.d_bresp(split15_merge15_bresp[1:0])
    ,.d_bvalid(split15_merge15_bvalid)
    ,.d_rdata(split15_merge15_rdata[(DWID - 1):0])
    ,.d_rid(split15_merge15_rid[(IDWID - 1):0])
    ,.d_rlast(split15_merge15_rlast)
    ,.d_rready(split15_merge15_rready)
    ,.d_rresp(split15_merge15_rresp[1:0])
    ,.d_rvalid(split15_merge15_rvalid)
    ,.d_wdata(split15_merge15_wdata[(DWID - 1):0])
    ,.d_wlast(split15_merge15_wlast)
    ,.d_wready(split15_merge15_wready)
    ,.d_wstrb(split15_merge15_wstrb[(WSTRB - 1):0])
    ,.d_wvalid(split15_merge15_wvalid)
);


axi_4_splitter split13 (
     .clk(clk) ,.rst_n(rst_n)

    ,.araddr(mst13_araddr[31:0])
    ,.arburst(mst13_arburst[1:0])
    ,.arextras(mst13_arextras[(EXTRAS - 1):0])
    ,.arid(mst13_arid[(IDWID - 1):0])
    ,.arlen(mst13_arlen[7:0])
    ,.arready(mst13_arready)
    ,.arvalid(mst13_arvalid)
    ,.awaddr(mst13_awaddr[31:0])
    ,.awburst(mst13_awburst[1:0])
    ,.awextras(mst13_awextras[(EXTRAS - 1):0])
    ,.awid(mst13_awid[3:0])
    ,.awlen(mst13_awlen[7:0])
    ,.awready(mst13_awready)
    ,.awvalid(mst13_awvalid)
    ,.bid(mst13_bid[(IDWID - 1):0])
    ,.bready(mst13_bready)
    ,.bresp(mst13_bresp[1:0])
    ,.bvalid(mst13_bvalid)
    ,.rdata(mst13_rdata[(DWID - 1):0])
    ,.rid(mst13_rid[(IDWID - 1):0])
    ,.rlast(mst13_rlast)
    ,.rready(mst13_rready)
    ,.rresp(mst13_rresp[1:0])
    ,.rvalid(mst13_rvalid)
    ,.wdata(mst13_wdata[(DWID - 1):0])
    ,.wlast(mst13_wlast)
    ,.wready(mst13_wready)
    ,.wstrb(mst13_wstrb[(WSTRB - 1):0])
    ,.wvalid(mst13_wvalid)

    ,.a_araddr(split13_merge12_araddr[31:0])
    ,.a_arburst(split13_merge12_arburst[1:0])
    ,.a_arextras(split13_merge12_arextras[(EXTRAS - 1):0])
    ,.a_arid(split13_merge12_arid[(IDWID - 1):0])
    ,.a_arlen(split13_merge12_arlen[7:0])
    ,.a_arready(split13_merge12_arready)
    ,.a_arvalid(split13_merge12_arvalid)
    ,.a_awaddr(split13_merge12_awaddr[31:0])
    ,.a_awburst(split13_merge12_awburst[1:0])
    ,.a_awextras(split13_merge12_awextras[(EXTRAS - 1):0])
    ,.a_awid(split13_merge12_awid[(IDWID - 1):0])
    ,.a_awlen(split13_merge12_awlen[7:0])
    ,.a_awready(split13_merge12_awready)
    ,.a_awvalid(split13_merge12_awvalid)
    ,.a_bid(split13_merge12_bid[(IDWID - 1):0])
    ,.a_bready(split13_merge12_bready)
    ,.a_bresp(split13_merge12_bresp[1:0])
    ,.a_bvalid(split13_merge12_bvalid)
    ,.a_rdata(split13_merge12_rdata[(DWID - 1):0])
    ,.a_rid(split13_merge12_rid[(IDWID - 1):0])
    ,.a_rlast(split13_merge12_rlast)
    ,.a_rready(split13_merge12_rready)
    ,.a_rresp(split13_merge12_rresp[1:0])
    ,.a_rvalid(split13_merge12_rvalid)
    ,.a_wdata(split13_merge12_wdata[(DWID - 1):0])
    ,.a_wlast(split13_merge12_wlast)
    ,.a_wready(split13_merge12_wready)
    ,.a_wstrb(split13_merge12_wstrb[(WSTRB - 1):0])
    ,.a_wvalid(split13_merge12_wvalid)
    ,.b_araddr(split13_merge13_araddr[31:0])
    ,.b_arburst(split13_merge13_arburst[1:0])
    ,.b_arextras(split13_merge13_arextras[(EXTRAS - 1):0])
    ,.b_arid(split13_merge13_arid[(IDWID - 1):0])
    ,.b_arlen(split13_merge13_arlen[7:0])
    ,.b_arready(split13_merge13_arready)
    ,.b_arvalid(split13_merge13_arvalid)
    ,.b_awaddr(split13_merge13_awaddr[31:0])
    ,.b_awburst(split13_merge13_awburst[1:0])
    ,.b_awextras(split13_merge13_awextras[(EXTRAS - 1):0])
    ,.b_awid(split13_merge13_awid[(IDWID - 1):0])
    ,.b_awlen(split13_merge13_awlen[7:0])
    ,.b_awready(split13_merge13_awready)
    ,.b_awvalid(split13_merge13_awvalid)
    ,.b_bid(split13_merge13_bid[(IDWID - 1):0])
    ,.b_bready(split13_merge13_bready)
    ,.b_bresp(split13_merge13_bresp[1:0])
    ,.b_bvalid(split13_merge13_bvalid)
    ,.b_rdata(split13_merge13_rdata[(DWID - 1):0])
    ,.b_rid(split13_merge13_rid[(IDWID - 1):0])
    ,.b_rlast(split13_merge13_rlast)
    ,.b_rready(split13_merge13_rready)
    ,.b_rresp(split13_merge13_rresp[1:0])
    ,.b_rvalid(split13_merge13_rvalid)
    ,.b_wdata(split13_merge13_wdata[(DWID - 1):0])
    ,.b_wlast(split13_merge13_wlast)
    ,.b_wready(split13_merge13_wready)
    ,.b_wstrb(split13_merge13_wstrb[(WSTRB - 1):0])
    ,.b_wvalid(split13_merge13_wvalid)
    ,.c_araddr(split13_merge14_araddr[31:0])
    ,.c_arburst(split13_merge14_arburst[1:0])
    ,.c_arextras(split13_merge14_arextras[(EXTRAS - 1):0])
    ,.c_arid(split13_merge14_arid[(IDWID - 1):0])
    ,.c_arlen(split13_merge14_arlen[7:0])
    ,.c_arready(split13_merge14_arready)
    ,.c_arvalid(split13_merge14_arvalid)
    ,.c_awaddr(split13_merge14_awaddr[31:0])
    ,.c_awburst(split13_merge14_awburst[1:0])
    ,.c_awextras(split13_merge14_awextras[(EXTRAS - 1):0])
    ,.c_awid(split13_merge14_awid[(IDWID - 1):0])
    ,.c_awlen(split13_merge14_awlen[7:0])
    ,.c_awready(split13_merge14_awready)
    ,.c_awvalid(split13_merge14_awvalid)
    ,.c_bid(split13_merge14_bid[(IDWID - 1):0])
    ,.c_bready(split13_merge14_bready)
    ,.c_bresp(split13_merge14_bresp[1:0])
    ,.c_bvalid(split13_merge14_bvalid)
    ,.c_rdata(split13_merge14_rdata[(DWID - 1):0])
    ,.c_rid(split13_merge14_rid[(IDWID - 1):0])
    ,.c_rlast(split13_merge14_rlast)
    ,.c_rready(split13_merge14_rready)
    ,.c_rresp(split13_merge14_rresp[1:0])
    ,.c_rvalid(split13_merge14_rvalid)
    ,.c_wdata(split13_merge14_wdata[(DWID - 1):0])
    ,.c_wlast(split13_merge14_wlast)
    ,.c_wready(split13_merge14_wready)
    ,.c_wstrb(split13_merge14_wstrb[(WSTRB - 1):0])
    ,.c_wvalid(split13_merge14_wvalid)
    ,.d_araddr(split13_merge15_araddr[31:0])
    ,.d_arburst(split13_merge15_arburst[1:0])
    ,.d_arextras(split13_merge15_arextras[(EXTRAS - 1):0])
    ,.d_arid(split13_merge15_arid[(IDWID - 1):0])
    ,.d_arlen(split13_merge15_arlen[7:0])
    ,.d_arready(split13_merge15_arready)
    ,.d_arvalid(split13_merge15_arvalid)
    ,.d_awaddr(split13_merge15_awaddr[31:0])
    ,.d_awburst(split13_merge15_awburst[1:0])
    ,.d_awextras(split13_merge15_awextras[(EXTRAS - 1):0])
    ,.d_awid(split13_merge15_awid[(IDWID - 1):0])
    ,.d_awlen(split13_merge15_awlen[7:0])
    ,.d_awready(split13_merge15_awready)
    ,.d_awvalid(split13_merge15_awvalid)
    ,.d_bid(split13_merge15_bid[(IDWID - 1):0])
    ,.d_bready(split13_merge15_bready)
    ,.d_bresp(split13_merge15_bresp[1:0])
    ,.d_bvalid(split13_merge15_bvalid)
    ,.d_rdata(split13_merge15_rdata[(DWID - 1):0])
    ,.d_rid(split13_merge15_rid[(IDWID - 1):0])
    ,.d_rlast(split13_merge15_rlast)
    ,.d_rready(split13_merge15_rready)
    ,.d_rresp(split13_merge15_rresp[1:0])
    ,.d_rvalid(split13_merge15_rvalid)
    ,.d_wdata(split13_merge15_wdata[(DWID - 1):0])
    ,.d_wlast(split13_merge15_wlast)
    ,.d_wready(split13_merge15_wready)
    ,.d_wstrb(split13_merge15_wstrb[(WSTRB - 1):0])
    ,.d_wvalid(split13_merge15_wvalid)

);

axi_4_splitter split14 (
     .clk(clk) ,.rst_n(rst_n)

    ,.araddr(mst14_araddr[31:0])
    ,.arburst(mst14_arburst[1:0])
    ,.arextras(mst14_arextras[(EXTRAS - 1):0])
    ,.arid(mst14_arid[(IDWID - 1):0])
    ,.arlen(mst14_arlen[7:0])
    ,.arready(mst14_arready)
    ,.arvalid(mst14_arvalid)
    ,.awaddr(mst14_awaddr[31:0])
    ,.awburst(mst14_awburst[1:0])
    ,.awextras(mst14_awextras[(EXTRAS - 1):0])
    ,.awid(mst14_awid[3:0])
    ,.awlen(mst14_awlen[7:0])
    ,.awready(mst14_awready)
    ,.awvalid(mst14_awvalid)
    ,.bid(mst14_bid[(IDWID - 1):0])
    ,.bready(mst14_bready)
    ,.bresp(mst14_bresp[1:0])
    ,.bvalid(mst14_bvalid)
    ,.rdata(mst14_rdata[(DWID - 1):0])
    ,.rid(mst14_rid[(IDWID - 1):0])
    ,.rlast(mst14_rlast)
    ,.rready(mst14_rready)
    ,.rresp(mst14_rresp[1:0])
    ,.rvalid(mst14_rvalid)
    ,.wdata(mst14_wdata[(DWID - 1):0])
    ,.wlast(mst14_wlast)
    ,.wready(mst14_wready)
    ,.wstrb(mst14_wstrb[(WSTRB - 1):0])
    ,.wvalid(mst14_wvalid)

    ,.a_araddr(split14_merge12_araddr[31:0])
    ,.a_arburst(split14_merge12_arburst[1:0])
    ,.a_arextras(split14_merge12_arextras[(EXTRAS - 1):0])
    ,.a_arid(split14_merge12_arid[(IDWID - 1):0])
    ,.a_arlen(split14_merge12_arlen[7:0])
    ,.a_arready(split14_merge12_arready)
    ,.a_arvalid(split14_merge12_arvalid)
    ,.a_awaddr(split14_merge12_awaddr[31:0])
    ,.a_awburst(split14_merge12_awburst[1:0])
    ,.a_awextras(split14_merge12_awextras[(EXTRAS - 1):0])
    ,.a_awid(split14_merge12_awid[(IDWID - 1):0])
    ,.a_awlen(split14_merge12_awlen[7:0])
    ,.a_awready(split14_merge12_awready)
    ,.a_awvalid(split14_merge12_awvalid)
    ,.a_bid(split14_merge12_bid[(IDWID - 1):0])
    ,.a_bready(split14_merge12_bready)
    ,.a_bresp(split14_merge12_bresp[1:0])
    ,.a_bvalid(split14_merge12_bvalid)
    ,.a_rdata(split14_merge12_rdata[(DWID - 1):0])
    ,.a_rid(split14_merge12_rid[(IDWID - 1):0])
    ,.a_rlast(split14_merge12_rlast)
    ,.a_rready(split14_merge12_rready)
    ,.a_rresp(split14_merge12_rresp[1:0])
    ,.a_rvalid(split14_merge12_rvalid)
    ,.a_wdata(split14_merge12_wdata[(DWID - 1):0])
    ,.a_wlast(split14_merge12_wlast)
    ,.a_wready(split14_merge12_wready)
    ,.a_wstrb(split14_merge12_wstrb[(WSTRB - 1):0])
    ,.a_wvalid(split14_merge12_wvalid)
    ,.b_araddr(split14_merge13_araddr[31:0])
    ,.b_arburst(split14_merge13_arburst[1:0])
    ,.b_arextras(split14_merge13_arextras[(EXTRAS - 1):0])
    ,.b_arid(split14_merge13_arid[(IDWID - 1):0])
    ,.b_arlen(split14_merge13_arlen[7:0])
    ,.b_arready(split14_merge13_arready)
    ,.b_arvalid(split14_merge13_arvalid)
    ,.b_awaddr(split14_merge13_awaddr[31:0])
    ,.b_awburst(split14_merge13_awburst[1:0])
    ,.b_awextras(split14_merge13_awextras[(EXTRAS - 1):0])
    ,.b_awid(split14_merge13_awid[(IDWID - 1):0])
    ,.b_awlen(split14_merge13_awlen[7:0])
    ,.b_awready(split14_merge13_awready)
    ,.b_awvalid(split14_merge13_awvalid)
    ,.b_bid(split14_merge13_bid[(IDWID - 1):0])
    ,.b_bready(split14_merge13_bready)
    ,.b_bresp(split14_merge13_bresp[1:0])
    ,.b_bvalid(split14_merge13_bvalid)
    ,.b_rdata(split14_merge13_rdata[(DWID - 1):0])
    ,.b_rid(split14_merge13_rid[(IDWID - 1):0])
    ,.b_rlast(split14_merge13_rlast)
    ,.b_rready(split14_merge13_rready)
    ,.b_rresp(split14_merge13_rresp[1:0])
    ,.b_rvalid(split14_merge13_rvalid)
    ,.b_wdata(split14_merge13_wdata[(DWID - 1):0])
    ,.b_wlast(split14_merge13_wlast)
    ,.b_wready(split14_merge13_wready)
    ,.b_wstrb(split14_merge13_wstrb[(WSTRB - 1):0])
    ,.b_wvalid(split14_merge13_wvalid)
    ,.c_araddr(split14_merge14_araddr[31:0])
    ,.c_arburst(split14_merge14_arburst[1:0])
    ,.c_arextras(split14_merge14_arextras[(EXTRAS - 1):0])
    ,.c_arid(split14_merge14_arid[(IDWID - 1):0])
    ,.c_arlen(split14_merge14_arlen[7:0])
    ,.c_arready(split14_merge14_arready)
    ,.c_arvalid(split14_merge14_arvalid)
    ,.c_awaddr(split14_merge14_awaddr[31:0])
    ,.c_awburst(split14_merge14_awburst[1:0])
    ,.c_awextras(split14_merge14_awextras[(EXTRAS - 1):0])
    ,.c_awid(split14_merge14_awid[(IDWID - 1):0])
    ,.c_awlen(split14_merge14_awlen[7:0])
    ,.c_awready(split14_merge14_awready)
    ,.c_awvalid(split14_merge14_awvalid)
    ,.c_bid(split14_merge14_bid[(IDWID - 1):0])
    ,.c_bready(split14_merge14_bready)
    ,.c_bresp(split14_merge14_bresp[1:0])
    ,.c_bvalid(split14_merge14_bvalid)
    ,.c_rdata(split14_merge14_rdata[(DWID - 1):0])
    ,.c_rid(split14_merge14_rid[(IDWID - 1):0])
    ,.c_rlast(split14_merge14_rlast)
    ,.c_rready(split14_merge14_rready)
    ,.c_rresp(split14_merge14_rresp[1:0])
    ,.c_rvalid(split14_merge14_rvalid)
    ,.c_wdata(split14_merge14_wdata[(DWID - 1):0])
    ,.c_wlast(split14_merge14_wlast)
    ,.c_wready(split14_merge14_wready)
    ,.c_wstrb(split14_merge14_wstrb[(WSTRB - 1):0])
    ,.c_wvalid(split14_merge14_wvalid)
    ,.d_araddr(split14_merge15_araddr[31:0])
    ,.d_arburst(split14_merge15_arburst[1:0])
    ,.d_arextras(split14_merge15_arextras[(EXTRAS - 1):0])
    ,.d_arid(split14_merge15_arid[(IDWID - 1):0])
    ,.d_arlen(split14_merge15_arlen[7:0])
    ,.d_arready(split14_merge15_arready)
    ,.d_arvalid(split14_merge15_arvalid)
    ,.d_awaddr(split14_merge15_awaddr[31:0])
    ,.d_awburst(split14_merge15_awburst[1:0])
    ,.d_awextras(split14_merge15_awextras[(EXTRAS - 1):0])
    ,.d_awid(split14_merge15_awid[(IDWID - 1):0])
    ,.d_awlen(split14_merge15_awlen[7:0])
    ,.d_awready(split14_merge15_awready)
    ,.d_awvalid(split14_merge15_awvalid)
    ,.d_bid(split14_merge15_bid[(IDWID - 1):0])
    ,.d_bready(split14_merge15_bready)
    ,.d_bresp(split14_merge15_bresp[1:0])
    ,.d_bvalid(split14_merge15_bvalid)
    ,.d_rdata(split14_merge15_rdata[(DWID - 1):0])
    ,.d_rid(split14_merge15_rid[(IDWID - 1):0])
    ,.d_rlast(split14_merge15_rlast)
    ,.d_rready(split14_merge15_rready)
    ,.d_rresp(split14_merge15_rresp[1:0])
    ,.d_rvalid(split14_merge15_rvalid)
    ,.d_wdata(split14_merge15_wdata[(DWID - 1):0])
    ,.d_wlast(split14_merge15_wlast)
    ,.d_wready(split14_merge15_wready)
    ,.d_wstrb(split14_merge15_wstrb[(WSTRB - 1):0])
    ,.d_wvalid(split14_merge15_wvalid)

);

axi_4_splitter split15 (
     .clk(clk) ,.rst_n(rst_n)

    ,.araddr(mst15_araddr[31:0])
    ,.arburst(mst15_arburst[1:0])
    ,.arextras(mst15_arextras[(EXTRAS - 1):0])
    ,.arid(mst15_arid[(IDWID - 1):0])
    ,.arlen(mst15_arlen[7:0])
    ,.arready(mst15_arready)
    ,.arvalid(mst15_arvalid)
    ,.awaddr(mst15_awaddr[31:0])
    ,.awburst(mst15_awburst[1:0])
    ,.awextras(mst15_awextras[(EXTRAS - 1):0])
    ,.awid(mst15_awid[3:0])
    ,.awlen(mst15_awlen[7:0])
    ,.awready(mst15_awready)
    ,.awvalid(mst15_awvalid)
    ,.bid(mst15_bid[(IDWID - 1):0])
    ,.bready(mst15_bready)
    ,.bresp(mst15_bresp[1:0])
    ,.bvalid(mst15_bvalid)
    ,.rdata(mst15_rdata[(DWID - 1):0])
    ,.rid(mst15_rid[(IDWID - 1):0])
    ,.rlast(mst15_rlast)
    ,.rready(mst15_rready)
    ,.rresp(mst15_rresp[1:0])
    ,.rvalid(mst15_rvalid)
    ,.wdata(mst15_wdata[(DWID - 1):0])
    ,.wlast(mst15_wlast)
    ,.wready(mst15_wready)
    ,.wstrb(mst15_wstrb[(WSTRB - 1):0])
    ,.wvalid(mst15_wvalid)

    ,.a_araddr(split15_merge12_araddr[31:0])
    ,.a_arburst(split15_merge12_arburst[1:0])
    ,.a_arextras(split15_merge12_arextras[(EXTRAS - 1):0])
    ,.a_arid(split15_merge12_arid[(IDWID - 1):0])
    ,.a_arlen(split15_merge12_arlen[7:0])
    ,.a_arready(split15_merge12_arready)
    ,.a_arvalid(split15_merge12_arvalid)
    ,.a_awaddr(split15_merge12_awaddr[31:0])
    ,.a_awburst(split15_merge12_awburst[1:0])
    ,.a_awextras(split15_merge12_awextras[(EXTRAS - 1):0])
    ,.a_awid(split15_merge12_awid[(IDWID - 1):0])
    ,.a_awlen(split15_merge12_awlen[7:0])
    ,.a_awready(split15_merge12_awready)
    ,.a_awvalid(split15_merge12_awvalid)
    ,.a_bid(split15_merge12_bid[(IDWID - 1):0])
    ,.a_bready(split15_merge12_bready)
    ,.a_bresp(split15_merge12_bresp[1:0])
    ,.a_bvalid(split15_merge12_bvalid)
    ,.a_rdata(split15_merge12_rdata[(DWID - 1):0])
    ,.a_rid(split15_merge12_rid[(IDWID - 1):0])
    ,.a_rlast(split15_merge12_rlast)
    ,.a_rready(split15_merge12_rready)
    ,.a_rresp(split15_merge12_rresp[1:0])
    ,.a_rvalid(split15_merge12_rvalid)
    ,.a_wdata(split15_merge12_wdata[(DWID - 1):0])
    ,.a_wlast(split15_merge12_wlast)
    ,.a_wready(split15_merge12_wready)
    ,.a_wstrb(split15_merge12_wstrb[(WSTRB - 1):0])
    ,.a_wvalid(split15_merge12_wvalid)
    ,.b_araddr(split15_merge13_araddr[31:0])
    ,.b_arburst(split15_merge13_arburst[1:0])
    ,.b_arextras(split15_merge13_arextras[(EXTRAS - 1):0])
    ,.b_arid(split15_merge13_arid[(IDWID - 1):0])
    ,.b_arlen(split15_merge13_arlen[7:0])
    ,.b_arready(split15_merge13_arready)
    ,.b_arvalid(split15_merge13_arvalid)
    ,.b_awaddr(split15_merge13_awaddr[31:0])
    ,.b_awburst(split15_merge13_awburst[1:0])
    ,.b_awextras(split15_merge13_awextras[(EXTRAS - 1):0])
    ,.b_awid(split15_merge13_awid[(IDWID - 1):0])
    ,.b_awlen(split15_merge13_awlen[7:0])
    ,.b_awready(split15_merge13_awready)
    ,.b_awvalid(split15_merge13_awvalid)
    ,.b_bid(split15_merge13_bid[(IDWID - 1):0])
    ,.b_bready(split15_merge13_bready)
    ,.b_bresp(split15_merge13_bresp[1:0])
    ,.b_bvalid(split15_merge13_bvalid)
    ,.b_rdata(split15_merge13_rdata[(DWID - 1):0])
    ,.b_rid(split15_merge13_rid[(IDWID - 1):0])
    ,.b_rlast(split15_merge13_rlast)
    ,.b_rready(split15_merge13_rready)
    ,.b_rresp(split15_merge13_rresp[1:0])
    ,.b_rvalid(split15_merge13_rvalid)
    ,.b_wdata(split15_merge13_wdata[(DWID - 1):0])
    ,.b_wlast(split15_merge13_wlast)
    ,.b_wready(split15_merge13_wready)
    ,.b_wstrb(split15_merge13_wstrb[(WSTRB - 1):0])
    ,.b_wvalid(split15_merge13_wvalid)
    ,.c_araddr(split15_merge14_araddr[31:0])
    ,.c_arburst(split15_merge14_arburst[1:0])
    ,.c_arextras(split15_merge14_arextras[(EXTRAS - 1):0])
    ,.c_arid(split15_merge14_arid[(IDWID - 1):0])
    ,.c_arlen(split15_merge14_arlen[7:0])
    ,.c_arready(split15_merge14_arready)
    ,.c_arvalid(split15_merge14_arvalid)
    ,.c_awaddr(split15_merge14_awaddr[31:0])
    ,.c_awburst(split15_merge14_awburst[1:0])
    ,.c_awextras(split15_merge14_awextras[(EXTRAS - 1):0])
    ,.c_awid(split15_merge14_awid[(IDWID - 1):0])
    ,.c_awlen(split15_merge14_awlen[7:0])
    ,.c_awready(split15_merge14_awready)
    ,.c_awvalid(split15_merge14_awvalid)
    ,.c_bid(split15_merge14_bid[(IDWID - 1):0])
    ,.c_bready(split15_merge14_bready)
    ,.c_bresp(split15_merge14_bresp[1:0])
    ,.c_bvalid(split15_merge14_bvalid)
    ,.c_rdata(split15_merge14_rdata[(DWID - 1):0])
    ,.c_rid(split15_merge14_rid[(IDWID - 1):0])
    ,.c_rlast(split15_merge14_rlast)
    ,.c_rready(split15_merge14_rready)
    ,.c_rresp(split15_merge14_rresp[1:0])
    ,.c_rvalid(split15_merge14_rvalid)
    ,.c_wdata(split15_merge14_wdata[(DWID - 1):0])
    ,.c_wlast(split15_merge14_wlast)
    ,.c_wready(split15_merge14_wready)
    ,.c_wstrb(split15_merge14_wstrb[(WSTRB - 1):0])
    ,.c_wvalid(split15_merge14_wvalid)
    ,.d_araddr(split15_merge15_araddr[31:0])
    ,.d_arburst(split15_merge15_arburst[1:0])
    ,.d_arextras(split15_merge15_arextras[(EXTRAS - 1):0])
    ,.d_arid(split15_merge15_arid[(IDWID - 1):0])
    ,.d_arlen(split15_merge15_arlen[7:0])
    ,.d_arready(split15_merge15_arready)
    ,.d_arvalid(split15_merge15_arvalid)
    ,.d_awaddr(split15_merge15_awaddr[31:0])
    ,.d_awburst(split15_merge15_awburst[1:0])
    ,.d_awextras(split15_merge15_awextras[(EXTRAS - 1):0])
    ,.d_awid(split15_merge15_awid[(IDWID - 1):0])
    ,.d_awlen(split15_merge15_awlen[7:0])
    ,.d_awready(split15_merge15_awready)
    ,.d_awvalid(split15_merge15_awvalid)
    ,.d_bid(split15_merge15_bid[(IDWID - 1):0])
    ,.d_bready(split15_merge15_bready)
    ,.d_bresp(split15_merge15_bresp[1:0])
    ,.d_bvalid(split15_merge15_bvalid)
    ,.d_rdata(split15_merge15_rdata[(DWID - 1):0])
    ,.d_rid(split15_merge15_rid[(IDWID - 1):0])
    ,.d_rlast(split15_merge15_rlast)
    ,.d_rready(split15_merge15_rready)
    ,.d_rresp(split15_merge15_rresp[1:0])
    ,.d_rvalid(split15_merge15_rvalid)
    ,.d_wdata(split15_merge15_wdata[(DWID - 1):0])
    ,.d_wlast(split15_merge15_wlast)
    ,.d_wready(split15_merge15_wready)
    ,.d_wstrb(split15_merge15_wstrb[(WSTRB - 1):0])
    ,.d_wvalid(split15_merge15_wvalid)

);

wire [IDWID-1:0] split100_merge208_arid ;
wire [31:0] split100_merge208_araddr ;
wire [7:0] split100_merge208_arlen ;
wire [EXTRAS-1:0] split100_merge208_arextras ;
wire [1:0] split100_merge208_arburst ;
wire split100_merge208_arvalid ;
wire split100_merge208_arready ;
wire [IDWID-1:0] split100_merge208_rid ;
wire [DWID-1:0] split100_merge208_rdata ;
wire [1:0] split100_merge208_rresp ;
wire split100_merge208_rlast ;
wire split100_merge208_rvalid ;
wire split100_merge208_rready ;

wire [IDWID-1:0] split100_merge208_awid ;
wire [31:0] split100_merge208_awaddr ;
wire [7:0] split100_merge208_awlen ;
wire [EXTRAS-1:0] split100_merge208_awextras ;
wire [1:0] split100_merge208_awburst ;
wire split100_merge208_awvalid ;
wire split100_merge208_awready ;
wire [DWID-1:0] split100_merge208_wdata ;
wire [WSTRB-1:0] split100_merge208_wstrb ;
wire split100_merge208_wlast ;
wire split100_merge208_wvalid ;
wire split100_merge208_wready ;
wire [IDWID-1:0] split100_merge208_bid ;
wire [1:0] split100_merge208_bresp ;
wire split100_merge208_bvalid ;
wire split100_merge208_bready ;


wire [IDWID-1:0] split100_merge211_arid ;
wire [31:0] split100_merge211_araddr ;
wire [7:0] split100_merge211_arlen ;
wire [EXTRAS-1:0] split100_merge211_arextras ;
wire [1:0] split100_merge211_arburst ;
wire split100_merge211_arvalid ;
wire split100_merge211_arready ;
wire [IDWID-1:0] split100_merge211_rid ;
wire [DWID-1:0] split100_merge211_rdata ;
wire [1:0] split100_merge211_rresp ;
wire split100_merge211_rlast ;
wire split100_merge211_rvalid ;
wire split100_merge211_rready ;

wire [IDWID-1:0] split100_merge211_awid ;
wire [31:0] split100_merge211_awaddr ;
wire [7:0] split100_merge211_awlen ;
wire [EXTRAS-1:0] split100_merge211_awextras ;
wire [1:0] split100_merge211_awburst ;
wire split100_merge211_awvalid ;
wire split100_merge211_awready ;
wire [DWID-1:0] split100_merge211_wdata ;
wire [WSTRB-1:0] split100_merge211_wstrb ;
wire split100_merge211_wlast ;
wire split100_merge211_wvalid ;
wire split100_merge211_wready ;
wire [IDWID-1:0] split100_merge211_bid ;
wire [1:0] split100_merge211_bresp ;
wire split100_merge211_bvalid ;
wire split100_merge211_bready ;


wire [IDWID-1:0] split100_merge212_arid ;
wire [31:0] split100_merge212_araddr ;
wire [7:0] split100_merge212_arlen ;
wire [EXTRAS-1:0] split100_merge212_arextras ;
wire [1:0] split100_merge212_arburst ;
wire split100_merge212_arvalid ;
wire split100_merge212_arready ;
wire [IDWID-1:0] split100_merge212_rid ;
wire [DWID-1:0] split100_merge212_rdata ;
wire [1:0] split100_merge212_rresp ;
wire split100_merge212_rlast ;
wire split100_merge212_rvalid ;
wire split100_merge212_rready ;

wire [IDWID-1:0] split100_merge212_awid ;
wire [31:0] split100_merge212_awaddr ;
wire [7:0] split100_merge212_awlen ;
wire [EXTRAS-1:0] split100_merge212_awextras ;
wire [1:0] split100_merge212_awburst ;
wire split100_merge212_awvalid ;
wire split100_merge212_awready ;
wire [DWID-1:0] split100_merge212_wdata ;
wire [WSTRB-1:0] split100_merge212_wstrb ;
wire split100_merge212_wlast ;
wire split100_merge212_wvalid ;
wire split100_merge212_wready ;
wire [IDWID-1:0] split100_merge212_bid ;
wire [1:0] split100_merge212_bresp ;
wire split100_merge212_bvalid ;
wire split100_merge212_bready ;


wire [IDWID-1:0] split100_merge206_arid ;
wire [31:0] split100_merge206_araddr ;
wire [7:0] split100_merge206_arlen ;
wire [EXTRAS-1:0] split100_merge206_arextras ;
wire [1:0] split100_merge206_arburst ;
wire split100_merge206_arvalid ;
wire split100_merge206_arready ;
wire [IDWID-1:0] split100_merge206_rid ;
wire [DWID-1:0] split100_merge206_rdata ;
wire [1:0] split100_merge206_rresp ;
wire split100_merge206_rlast ;
wire split100_merge206_rvalid ;
wire split100_merge206_rready ;

wire [IDWID-1:0] split100_merge206_awid ;
wire [31:0] split100_merge206_awaddr ;
wire [7:0] split100_merge206_awlen ;
wire [EXTRAS-1:0] split100_merge206_awextras ;
wire [1:0] split100_merge206_awburst ;
wire split100_merge206_awvalid ;
wire split100_merge206_awready ;
wire [DWID-1:0] split100_merge206_wdata ;
wire [WSTRB-1:0] split100_merge206_wstrb ;
wire split100_merge206_wlast ;
wire split100_merge206_wvalid ;
wire split100_merge206_wready ;
wire [IDWID-1:0] split100_merge206_bid ;
wire [1:0] split100_merge206_bresp ;
wire split100_merge206_bvalid ;
wire split100_merge206_bready ;


axi_4_splitter split100 (
     .clk(clk) ,.rst_n(rst_n)

    ,.araddr(merge0_split100_araddr[31:0])
    ,.arburst(merge0_split100_arburst[1:0])
    ,.arextras(merge0_split100_arextras[(EXTRAS - 1):0])
    ,.arid(merge0_split100_arid[(IDWID - 1):0])
    ,.arlen(merge0_split100_arlen[7:0])
    ,.arready(merge0_split100_arready)
    ,.arvalid(merge0_split100_arvalid)
    ,.awaddr(merge0_split100_awaddr[31:0])
    ,.awburst(merge0_split100_awburst[1:0])
    ,.awextras(merge0_split100_awextras[(EXTRAS - 1):0])
    ,.awid(merge0_split100_awid[3:0])
    ,.awlen(merge0_split100_awlen[7:0])
    ,.awready(merge0_split100_awready)
    ,.awvalid(merge0_split100_awvalid)
    ,.bid(merge0_split100_bid[(IDWID - 1):0])
    ,.bready(merge0_split100_bready)
    ,.bresp(merge0_split100_bresp[1:0])
    ,.bvalid(merge0_split100_bvalid)
    ,.rdata(merge0_split100_rdata[(DWID - 1):0])
    ,.rid(merge0_split100_rid[(IDWID - 1):0])
    ,.rlast(merge0_split100_rlast)
    ,.rready(merge0_split100_rready)
    ,.rresp(merge0_split100_rresp[1:0])
    ,.rvalid(merge0_split100_rvalid)
    ,.wdata(merge0_split100_wdata[(DWID - 1):0])
    ,.wlast(merge0_split100_wlast)
    ,.wready(merge0_split100_wready)
    ,.wstrb(merge0_split100_wstrb[(WSTRB - 1):0])
    ,.wvalid(merge0_split100_wvalid)

    ,.a_araddr(split100_merge208_araddr[31:0])
    ,.a_arburst(split100_merge208_arburst[1:0])
    ,.a_arextras(split100_merge208_arextras[(EXTRAS - 1):0])
    ,.a_arid(split100_merge208_arid[(IDWID - 1):0])
    ,.a_arlen(split100_merge208_arlen[7:0])
    ,.a_arready(split100_merge208_arready)
    ,.a_arvalid(split100_merge208_arvalid)
    ,.a_awaddr(split100_merge208_awaddr[31:0])
    ,.a_awburst(split100_merge208_awburst[1:0])
    ,.a_awextras(split100_merge208_awextras[(EXTRAS - 1):0])
    ,.a_awid(split100_merge208_awid[(IDWID - 1):0])
    ,.a_awlen(split100_merge208_awlen[7:0])
    ,.a_awready(split100_merge208_awready)
    ,.a_awvalid(split100_merge208_awvalid)
    ,.a_bid(split100_merge208_bid[(IDWID - 1):0])
    ,.a_bready(split100_merge208_bready)
    ,.a_bresp(split100_merge208_bresp[1:0])
    ,.a_bvalid(split100_merge208_bvalid)
    ,.a_rdata(split100_merge208_rdata[(DWID - 1):0])
    ,.a_rid(split100_merge208_rid[(IDWID - 1):0])
    ,.a_rlast(split100_merge208_rlast)
    ,.a_rready(split100_merge208_rready)
    ,.a_rresp(split100_merge208_rresp[1:0])
    ,.a_rvalid(split100_merge208_rvalid)
    ,.a_wdata(split100_merge208_wdata[(DWID - 1):0])
    ,.a_wlast(split100_merge208_wlast)
    ,.a_wready(split100_merge208_wready)
    ,.a_wstrb(split100_merge208_wstrb[(WSTRB - 1):0])
    ,.a_wvalid(split100_merge208_wvalid)
    ,.b_araddr(split100_merge211_araddr[31:0])
    ,.b_arburst(split100_merge211_arburst[1:0])
    ,.b_arextras(split100_merge211_arextras[(EXTRAS - 1):0])
    ,.b_arid(split100_merge211_arid[(IDWID - 1):0])
    ,.b_arlen(split100_merge211_arlen[7:0])
    ,.b_arready(split100_merge211_arready)
    ,.b_arvalid(split100_merge211_arvalid)
    ,.b_awaddr(split100_merge211_awaddr[31:0])
    ,.b_awburst(split100_merge211_awburst[1:0])
    ,.b_awextras(split100_merge211_awextras[(EXTRAS - 1):0])
    ,.b_awid(split100_merge211_awid[(IDWID - 1):0])
    ,.b_awlen(split100_merge211_awlen[7:0])
    ,.b_awready(split100_merge211_awready)
    ,.b_awvalid(split100_merge211_awvalid)
    ,.b_bid(split100_merge211_bid[(IDWID - 1):0])
    ,.b_bready(split100_merge211_bready)
    ,.b_bresp(split100_merge211_bresp[1:0])
    ,.b_bvalid(split100_merge211_bvalid)
    ,.b_rdata(split100_merge211_rdata[(DWID - 1):0])
    ,.b_rid(split100_merge211_rid[(IDWID - 1):0])
    ,.b_rlast(split100_merge211_rlast)
    ,.b_rready(split100_merge211_rready)
    ,.b_rresp(split100_merge211_rresp[1:0])
    ,.b_rvalid(split100_merge211_rvalid)
    ,.b_wdata(split100_merge211_wdata[(DWID - 1):0])
    ,.b_wlast(split100_merge211_wlast)
    ,.b_wready(split100_merge211_wready)
    ,.b_wstrb(split100_merge211_wstrb[(WSTRB - 1):0])
    ,.b_wvalid(split100_merge211_wvalid)
    ,.c_araddr(split100_merge212_araddr[31:0])
    ,.c_arburst(split100_merge212_arburst[1:0])
    ,.c_arextras(split100_merge212_arextras[(EXTRAS - 1):0])
    ,.c_arid(split100_merge212_arid[(IDWID - 1):0])
    ,.c_arlen(split100_merge212_arlen[7:0])
    ,.c_arready(split100_merge212_arready)
    ,.c_arvalid(split100_merge212_arvalid)
    ,.c_awaddr(split100_merge212_awaddr[31:0])
    ,.c_awburst(split100_merge212_awburst[1:0])
    ,.c_awextras(split100_merge212_awextras[(EXTRAS - 1):0])
    ,.c_awid(split100_merge212_awid[(IDWID - 1):0])
    ,.c_awlen(split100_merge212_awlen[7:0])
    ,.c_awready(split100_merge212_awready)
    ,.c_awvalid(split100_merge212_awvalid)
    ,.c_bid(split100_merge212_bid[(IDWID - 1):0])
    ,.c_bready(split100_merge212_bready)
    ,.c_bresp(split100_merge212_bresp[1:0])
    ,.c_bvalid(split100_merge212_bvalid)
    ,.c_rdata(split100_merge212_rdata[(DWID - 1):0])
    ,.c_rid(split100_merge212_rid[(IDWID - 1):0])
    ,.c_rlast(split100_merge212_rlast)
    ,.c_rready(split100_merge212_rready)
    ,.c_rresp(split100_merge212_rresp[1:0])
    ,.c_rvalid(split100_merge212_rvalid)
    ,.c_wdata(split100_merge212_wdata[(DWID - 1):0])
    ,.c_wlast(split100_merge212_wlast)
    ,.c_wready(split100_merge212_wready)
    ,.c_wstrb(split100_merge212_wstrb[(WSTRB - 1):0])
    ,.c_wvalid(split100_merge212_wvalid)
    ,.d_araddr(split100_merge206_araddr[31:0])
    ,.d_arburst(split100_merge206_arburst[1:0])
    ,.d_arextras(split100_merge206_arextras[(EXTRAS - 1):0])
    ,.d_arid(split100_merge206_arid[(IDWID - 1):0])
    ,.d_arlen(split100_merge206_arlen[7:0])
    ,.d_arready(split100_merge206_arready)
    ,.d_arvalid(split100_merge206_arvalid)
    ,.d_awaddr(split100_merge206_awaddr[31:0])
    ,.d_awburst(split100_merge206_awburst[1:0])
    ,.d_awextras(split100_merge206_awextras[(EXTRAS - 1):0])
    ,.d_awid(split100_merge206_awid[(IDWID - 1):0])
    ,.d_awlen(split100_merge206_awlen[7:0])
    ,.d_awready(split100_merge206_awready)
    ,.d_awvalid(split100_merge206_awvalid)
    ,.d_bid(split100_merge206_bid[(IDWID - 1):0])
    ,.d_bready(split100_merge206_bready)
    ,.d_bresp(split100_merge206_bresp[1:0])
    ,.d_bvalid(split100_merge206_bvalid)
    ,.d_rdata(split100_merge206_rdata[(DWID - 1):0])
    ,.d_rid(split100_merge206_rid[(IDWID - 1):0])
    ,.d_rlast(split100_merge206_rlast)
    ,.d_rready(split100_merge206_rready)
    ,.d_rresp(split100_merge206_rresp[1:0])
    ,.d_rvalid(split100_merge206_rvalid)
    ,.d_wdata(split100_merge206_wdata[(DWID - 1):0])
    ,.d_wlast(split100_merge206_wlast)
    ,.d_wready(split100_merge206_wready)
    ,.d_wstrb(split100_merge206_wstrb[(WSTRB - 1):0])
    ,.d_wvalid(split100_merge206_wvalid)

);

wire [IDWID-1:0] split101_merge203_arid ;
wire [31:0] split101_merge203_araddr ;
wire [7:0] split101_merge203_arlen ;
wire [EXTRAS-1:0] split101_merge203_arextras ;
wire [1:0] split101_merge203_arburst ;
wire split101_merge203_arvalid ;
wire split101_merge203_arready ;
wire [IDWID-1:0] split101_merge203_rid ;
wire [DWID-1:0] split101_merge203_rdata ;
wire [1:0] split101_merge203_rresp ;
wire split101_merge203_rlast ;
wire split101_merge203_rvalid ;
wire split101_merge203_rready ;

wire [IDWID-1:0] split101_merge203_awid ;
wire [31:0] split101_merge203_awaddr ;
wire [7:0] split101_merge203_awlen ;
wire [EXTRAS-1:0] split101_merge203_awextras ;
wire [1:0] split101_merge203_awburst ;
wire split101_merge203_awvalid ;
wire split101_merge203_awready ;
wire [DWID-1:0] split101_merge203_wdata ;
wire [WSTRB-1:0] split101_merge203_wstrb ;
wire split101_merge203_wlast ;
wire split101_merge203_wvalid ;
wire split101_merge203_wready ;
wire [IDWID-1:0] split101_merge203_bid ;
wire [1:0] split101_merge203_bresp ;
wire split101_merge203_bvalid ;
wire split101_merge203_bready ;


wire [IDWID-1:0] split101_merge201_arid ;
wire [31:0] split101_merge201_araddr ;
wire [7:0] split101_merge201_arlen ;
wire [EXTRAS-1:0] split101_merge201_arextras ;
wire [1:0] split101_merge201_arburst ;
wire split101_merge201_arvalid ;
wire split101_merge201_arready ;
wire [IDWID-1:0] split101_merge201_rid ;
wire [DWID-1:0] split101_merge201_rdata ;
wire [1:0] split101_merge201_rresp ;
wire split101_merge201_rlast ;
wire split101_merge201_rvalid ;
wire split101_merge201_rready ;

wire [IDWID-1:0] split101_merge201_awid ;
wire [31:0] split101_merge201_awaddr ;
wire [7:0] split101_merge201_awlen ;
wire [EXTRAS-1:0] split101_merge201_awextras ;
wire [1:0] split101_merge201_awburst ;
wire split101_merge201_awvalid ;
wire split101_merge201_awready ;
wire [DWID-1:0] split101_merge201_wdata ;
wire [WSTRB-1:0] split101_merge201_wstrb ;
wire split101_merge201_wlast ;
wire split101_merge201_wvalid ;
wire split101_merge201_wready ;
wire [IDWID-1:0] split101_merge201_bid ;
wire [1:0] split101_merge201_bresp ;
wire split101_merge201_bvalid ;
wire split101_merge201_bready ;


wire [IDWID-1:0] split101_merge212_arid ;
wire [31:0] split101_merge212_araddr ;
wire [7:0] split101_merge212_arlen ;
wire [EXTRAS-1:0] split101_merge212_arextras ;
wire [1:0] split101_merge212_arburst ;
wire split101_merge212_arvalid ;
wire split101_merge212_arready ;
wire [IDWID-1:0] split101_merge212_rid ;
wire [DWID-1:0] split101_merge212_rdata ;
wire [1:0] split101_merge212_rresp ;
wire split101_merge212_rlast ;
wire split101_merge212_rvalid ;
wire split101_merge212_rready ;

wire [IDWID-1:0] split101_merge212_awid ;
wire [31:0] split101_merge212_awaddr ;
wire [7:0] split101_merge212_awlen ;
wire [EXTRAS-1:0] split101_merge212_awextras ;
wire [1:0] split101_merge212_awburst ;
wire split101_merge212_awvalid ;
wire split101_merge212_awready ;
wire [DWID-1:0] split101_merge212_wdata ;
wire [WSTRB-1:0] split101_merge212_wstrb ;
wire split101_merge212_wlast ;
wire split101_merge212_wvalid ;
wire split101_merge212_wready ;
wire [IDWID-1:0] split101_merge212_bid ;
wire [1:0] split101_merge212_bresp ;
wire split101_merge212_bvalid ;
wire split101_merge212_bready ;


wire [IDWID-1:0] split101_merge209_arid ;
wire [31:0] split101_merge209_araddr ;
wire [7:0] split101_merge209_arlen ;
wire [EXTRAS-1:0] split101_merge209_arextras ;
wire [1:0] split101_merge209_arburst ;
wire split101_merge209_arvalid ;
wire split101_merge209_arready ;
wire [IDWID-1:0] split101_merge209_rid ;
wire [DWID-1:0] split101_merge209_rdata ;
wire [1:0] split101_merge209_rresp ;
wire split101_merge209_rlast ;
wire split101_merge209_rvalid ;
wire split101_merge209_rready ;

wire [IDWID-1:0] split101_merge209_awid ;
wire [31:0] split101_merge209_awaddr ;
wire [7:0] split101_merge209_awlen ;
wire [EXTRAS-1:0] split101_merge209_awextras ;
wire [1:0] split101_merge209_awburst ;
wire split101_merge209_awvalid ;
wire split101_merge209_awready ;
wire [DWID-1:0] split101_merge209_wdata ;
wire [WSTRB-1:0] split101_merge209_wstrb ;
wire split101_merge209_wlast ;
wire split101_merge209_wvalid ;
wire split101_merge209_wready ;
wire [IDWID-1:0] split101_merge209_bid ;
wire [1:0] split101_merge209_bresp ;
wire split101_merge209_bvalid ;
wire split101_merge209_bready ;


axi_4_splitter split101 (
     .clk(clk) ,.rst_n(rst_n)

    ,.araddr(merge1_split101_araddr[31:0])
    ,.arburst(merge1_split101_arburst[1:0])
    ,.arextras(merge1_split101_arextras[(EXTRAS - 1):0])
    ,.arid(merge1_split101_arid[(IDWID - 1):0])
    ,.arlen(merge1_split101_arlen[7:0])
    ,.arready(merge1_split101_arready)
    ,.arvalid(merge1_split101_arvalid)
    ,.awaddr(merge1_split101_awaddr[31:0])
    ,.awburst(merge1_split101_awburst[1:0])
    ,.awextras(merge1_split101_awextras[(EXTRAS - 1):0])
    ,.awid(merge1_split101_awid[3:0])
    ,.awlen(merge1_split101_awlen[7:0])
    ,.awready(merge1_split101_awready)
    ,.awvalid(merge1_split101_awvalid)
    ,.bid(merge1_split101_bid[(IDWID - 1):0])
    ,.bready(merge1_split101_bready)
    ,.bresp(merge1_split101_bresp[1:0])
    ,.bvalid(merge1_split101_bvalid)
    ,.rdata(merge1_split101_rdata[(DWID - 1):0])
    ,.rid(merge1_split101_rid[(IDWID - 1):0])
    ,.rlast(merge1_split101_rlast)
    ,.rready(merge1_split101_rready)
    ,.rresp(merge1_split101_rresp[1:0])
    ,.rvalid(merge1_split101_rvalid)
    ,.wdata(merge1_split101_wdata[(DWID - 1):0])
    ,.wlast(merge1_split101_wlast)
    ,.wready(merge1_split101_wready)
    ,.wstrb(merge1_split101_wstrb[(WSTRB - 1):0])
    ,.wvalid(merge1_split101_wvalid)

    ,.a_araddr(split101_merge203_araddr[31:0])
    ,.a_arburst(split101_merge203_arburst[1:0])
    ,.a_arextras(split101_merge203_arextras[(EXTRAS - 1):0])
    ,.a_arid(split101_merge203_arid[(IDWID - 1):0])
    ,.a_arlen(split101_merge203_arlen[7:0])
    ,.a_arready(split101_merge203_arready)
    ,.a_arvalid(split101_merge203_arvalid)
    ,.a_awaddr(split101_merge203_awaddr[31:0])
    ,.a_awburst(split101_merge203_awburst[1:0])
    ,.a_awextras(split101_merge203_awextras[(EXTRAS - 1):0])
    ,.a_awid(split101_merge203_awid[(IDWID - 1):0])
    ,.a_awlen(split101_merge203_awlen[7:0])
    ,.a_awready(split101_merge203_awready)
    ,.a_awvalid(split101_merge203_awvalid)
    ,.a_bid(split101_merge203_bid[(IDWID - 1):0])
    ,.a_bready(split101_merge203_bready)
    ,.a_bresp(split101_merge203_bresp[1:0])
    ,.a_bvalid(split101_merge203_bvalid)
    ,.a_rdata(split101_merge203_rdata[(DWID - 1):0])
    ,.a_rid(split101_merge203_rid[(IDWID - 1):0])
    ,.a_rlast(split101_merge203_rlast)
    ,.a_rready(split101_merge203_rready)
    ,.a_rresp(split101_merge203_rresp[1:0])
    ,.a_rvalid(split101_merge203_rvalid)
    ,.a_wdata(split101_merge203_wdata[(DWID - 1):0])
    ,.a_wlast(split101_merge203_wlast)
    ,.a_wready(split101_merge203_wready)
    ,.a_wstrb(split101_merge203_wstrb[(WSTRB - 1):0])
    ,.a_wvalid(split101_merge203_wvalid)
    ,.b_araddr(split101_merge201_araddr[31:0])
    ,.b_arburst(split101_merge201_arburst[1:0])
    ,.b_arextras(split101_merge201_arextras[(EXTRAS - 1):0])
    ,.b_arid(split101_merge201_arid[(IDWID - 1):0])
    ,.b_arlen(split101_merge201_arlen[7:0])
    ,.b_arready(split101_merge201_arready)
    ,.b_arvalid(split101_merge201_arvalid)
    ,.b_awaddr(split101_merge201_awaddr[31:0])
    ,.b_awburst(split101_merge201_awburst[1:0])
    ,.b_awextras(split101_merge201_awextras[(EXTRAS - 1):0])
    ,.b_awid(split101_merge201_awid[(IDWID - 1):0])
    ,.b_awlen(split101_merge201_awlen[7:0])
    ,.b_awready(split101_merge201_awready)
    ,.b_awvalid(split101_merge201_awvalid)
    ,.b_bid(split101_merge201_bid[(IDWID - 1):0])
    ,.b_bready(split101_merge201_bready)
    ,.b_bresp(split101_merge201_bresp[1:0])
    ,.b_bvalid(split101_merge201_bvalid)
    ,.b_rdata(split101_merge201_rdata[(DWID - 1):0])
    ,.b_rid(split101_merge201_rid[(IDWID - 1):0])
    ,.b_rlast(split101_merge201_rlast)
    ,.b_rready(split101_merge201_rready)
    ,.b_rresp(split101_merge201_rresp[1:0])
    ,.b_rvalid(split101_merge201_rvalid)
    ,.b_wdata(split101_merge201_wdata[(DWID - 1):0])
    ,.b_wlast(split101_merge201_wlast)
    ,.b_wready(split101_merge201_wready)
    ,.b_wstrb(split101_merge201_wstrb[(WSTRB - 1):0])
    ,.b_wvalid(split101_merge201_wvalid)
    ,.c_araddr(split101_merge212_araddr[31:0])
    ,.c_arburst(split101_merge212_arburst[1:0])
    ,.c_arextras(split101_merge212_arextras[(EXTRAS - 1):0])
    ,.c_arid(split101_merge212_arid[(IDWID - 1):0])
    ,.c_arlen(split101_merge212_arlen[7:0])
    ,.c_arready(split101_merge212_arready)
    ,.c_arvalid(split101_merge212_arvalid)
    ,.c_awaddr(split101_merge212_awaddr[31:0])
    ,.c_awburst(split101_merge212_awburst[1:0])
    ,.c_awextras(split101_merge212_awextras[(EXTRAS - 1):0])
    ,.c_awid(split101_merge212_awid[(IDWID - 1):0])
    ,.c_awlen(split101_merge212_awlen[7:0])
    ,.c_awready(split101_merge212_awready)
    ,.c_awvalid(split101_merge212_awvalid)
    ,.c_bid(split101_merge212_bid[(IDWID - 1):0])
    ,.c_bready(split101_merge212_bready)
    ,.c_bresp(split101_merge212_bresp[1:0])
    ,.c_bvalid(split101_merge212_bvalid)
    ,.c_rdata(split101_merge212_rdata[(DWID - 1):0])
    ,.c_rid(split101_merge212_rid[(IDWID - 1):0])
    ,.c_rlast(split101_merge212_rlast)
    ,.c_rready(split101_merge212_rready)
    ,.c_rresp(split101_merge212_rresp[1:0])
    ,.c_rvalid(split101_merge212_rvalid)
    ,.c_wdata(split101_merge212_wdata[(DWID - 1):0])
    ,.c_wlast(split101_merge212_wlast)
    ,.c_wready(split101_merge212_wready)
    ,.c_wstrb(split101_merge212_wstrb[(WSTRB - 1):0])
    ,.c_wvalid(split101_merge212_wvalid)
    ,.d_araddr(split101_merge209_araddr[31:0])
    ,.d_arburst(split101_merge209_arburst[1:0])
    ,.d_arextras(split101_merge209_arextras[(EXTRAS - 1):0])
    ,.d_arid(split101_merge209_arid[(IDWID - 1):0])
    ,.d_arlen(split101_merge209_arlen[7:0])
    ,.d_arready(split101_merge209_arready)
    ,.d_arvalid(split101_merge209_arvalid)
    ,.d_awaddr(split101_merge209_awaddr[31:0])
    ,.d_awburst(split101_merge209_awburst[1:0])
    ,.d_awextras(split101_merge209_awextras[(EXTRAS - 1):0])
    ,.d_awid(split101_merge209_awid[(IDWID - 1):0])
    ,.d_awlen(split101_merge209_awlen[7:0])
    ,.d_awready(split101_merge209_awready)
    ,.d_awvalid(split101_merge209_awvalid)
    ,.d_bid(split101_merge209_bid[(IDWID - 1):0])
    ,.d_bready(split101_merge209_bready)
    ,.d_bresp(split101_merge209_bresp[1:0])
    ,.d_bvalid(split101_merge209_bvalid)
    ,.d_rdata(split101_merge209_rdata[(DWID - 1):0])
    ,.d_rid(split101_merge209_rid[(IDWID - 1):0])
    ,.d_rlast(split101_merge209_rlast)
    ,.d_rready(split101_merge209_rready)
    ,.d_rresp(split101_merge209_rresp[1:0])
    ,.d_rvalid(split101_merge209_rvalid)
    ,.d_wdata(split101_merge209_wdata[(DWID - 1):0])
    ,.d_wlast(split101_merge209_wlast)
    ,.d_wready(split101_merge209_wready)
    ,.d_wstrb(split101_merge209_wstrb[(WSTRB - 1):0])
    ,.d_wvalid(split101_merge209_wvalid)

);

wire [IDWID-1:0] split102_merge201_arid ;
wire [31:0] split102_merge201_araddr ;
wire [7:0] split102_merge201_arlen ;
wire [EXTRAS-1:0] split102_merge201_arextras ;
wire [1:0] split102_merge201_arburst ;
wire split102_merge201_arvalid ;
wire split102_merge201_arready ;
wire [IDWID-1:0] split102_merge201_rid ;
wire [DWID-1:0] split102_merge201_rdata ;
wire [1:0] split102_merge201_rresp ;
wire split102_merge201_rlast ;
wire split102_merge201_rvalid ;
wire split102_merge201_rready ;

wire [IDWID-1:0] split102_merge201_awid ;
wire [31:0] split102_merge201_awaddr ;
wire [7:0] split102_merge201_awlen ;
wire [EXTRAS-1:0] split102_merge201_awextras ;
wire [1:0] split102_merge201_awburst ;
wire split102_merge201_awvalid ;
wire split102_merge201_awready ;
wire [DWID-1:0] split102_merge201_wdata ;
wire [WSTRB-1:0] split102_merge201_wstrb ;
wire split102_merge201_wlast ;
wire split102_merge201_wvalid ;
wire split102_merge201_wready ;
wire [IDWID-1:0] split102_merge201_bid ;
wire [1:0] split102_merge201_bresp ;
wire split102_merge201_bvalid ;
wire split102_merge201_bready ;


wire [IDWID-1:0] split102_merge200_arid ;
wire [31:0] split102_merge200_araddr ;
wire [7:0] split102_merge200_arlen ;
wire [EXTRAS-1:0] split102_merge200_arextras ;
wire [1:0] split102_merge200_arburst ;
wire split102_merge200_arvalid ;
wire split102_merge200_arready ;
wire [IDWID-1:0] split102_merge200_rid ;
wire [DWID-1:0] split102_merge200_rdata ;
wire [1:0] split102_merge200_rresp ;
wire split102_merge200_rlast ;
wire split102_merge200_rvalid ;
wire split102_merge200_rready ;

wire [IDWID-1:0] split102_merge200_awid ;
wire [31:0] split102_merge200_awaddr ;
wire [7:0] split102_merge200_awlen ;
wire [EXTRAS-1:0] split102_merge200_awextras ;
wire [1:0] split102_merge200_awburst ;
wire split102_merge200_awvalid ;
wire split102_merge200_awready ;
wire [DWID-1:0] split102_merge200_wdata ;
wire [WSTRB-1:0] split102_merge200_wstrb ;
wire split102_merge200_wlast ;
wire split102_merge200_wvalid ;
wire split102_merge200_wready ;
wire [IDWID-1:0] split102_merge200_bid ;
wire [1:0] split102_merge200_bresp ;
wire split102_merge200_bvalid ;
wire split102_merge200_bready ;


wire [IDWID-1:0] split102_merge207_arid ;
wire [31:0] split102_merge207_araddr ;
wire [7:0] split102_merge207_arlen ;
wire [EXTRAS-1:0] split102_merge207_arextras ;
wire [1:0] split102_merge207_arburst ;
wire split102_merge207_arvalid ;
wire split102_merge207_arready ;
wire [IDWID-1:0] split102_merge207_rid ;
wire [DWID-1:0] split102_merge207_rdata ;
wire [1:0] split102_merge207_rresp ;
wire split102_merge207_rlast ;
wire split102_merge207_rvalid ;
wire split102_merge207_rready ;

wire [IDWID-1:0] split102_merge207_awid ;
wire [31:0] split102_merge207_awaddr ;
wire [7:0] split102_merge207_awlen ;
wire [EXTRAS-1:0] split102_merge207_awextras ;
wire [1:0] split102_merge207_awburst ;
wire split102_merge207_awvalid ;
wire split102_merge207_awready ;
wire [DWID-1:0] split102_merge207_wdata ;
wire [WSTRB-1:0] split102_merge207_wstrb ;
wire split102_merge207_wlast ;
wire split102_merge207_wvalid ;
wire split102_merge207_wready ;
wire [IDWID-1:0] split102_merge207_bid ;
wire [1:0] split102_merge207_bresp ;
wire split102_merge207_bvalid ;
wire split102_merge207_bready ;


wire [IDWID-1:0] split102_merge205_arid ;
wire [31:0] split102_merge205_araddr ;
wire [7:0] split102_merge205_arlen ;
wire [EXTRAS-1:0] split102_merge205_arextras ;
wire [1:0] split102_merge205_arburst ;
wire split102_merge205_arvalid ;
wire split102_merge205_arready ;
wire [IDWID-1:0] split102_merge205_rid ;
wire [DWID-1:0] split102_merge205_rdata ;
wire [1:0] split102_merge205_rresp ;
wire split102_merge205_rlast ;
wire split102_merge205_rvalid ;
wire split102_merge205_rready ;

wire [IDWID-1:0] split102_merge205_awid ;
wire [31:0] split102_merge205_awaddr ;
wire [7:0] split102_merge205_awlen ;
wire [EXTRAS-1:0] split102_merge205_awextras ;
wire [1:0] split102_merge205_awburst ;
wire split102_merge205_awvalid ;
wire split102_merge205_awready ;
wire [DWID-1:0] split102_merge205_wdata ;
wire [WSTRB-1:0] split102_merge205_wstrb ;
wire split102_merge205_wlast ;
wire split102_merge205_wvalid ;
wire split102_merge205_wready ;
wire [IDWID-1:0] split102_merge205_bid ;
wire [1:0] split102_merge205_bresp ;
wire split102_merge205_bvalid ;
wire split102_merge205_bready ;


axi_4_splitter split102 (
     .clk(clk) ,.rst_n(rst_n)

    ,.araddr(merge2_split102_araddr[31:0])
    ,.arburst(merge2_split102_arburst[1:0])
    ,.arextras(merge2_split102_arextras[(EXTRAS - 1):0])
    ,.arid(merge2_split102_arid[(IDWID - 1):0])
    ,.arlen(merge2_split102_arlen[7:0])
    ,.arready(merge2_split102_arready)
    ,.arvalid(merge2_split102_arvalid)
    ,.awaddr(merge2_split102_awaddr[31:0])
    ,.awburst(merge2_split102_awburst[1:0])
    ,.awextras(merge2_split102_awextras[(EXTRAS - 1):0])
    ,.awid(merge2_split102_awid[3:0])
    ,.awlen(merge2_split102_awlen[7:0])
    ,.awready(merge2_split102_awready)
    ,.awvalid(merge2_split102_awvalid)
    ,.bid(merge2_split102_bid[(IDWID - 1):0])
    ,.bready(merge2_split102_bready)
    ,.bresp(merge2_split102_bresp[1:0])
    ,.bvalid(merge2_split102_bvalid)
    ,.rdata(merge2_split102_rdata[(DWID - 1):0])
    ,.rid(merge2_split102_rid[(IDWID - 1):0])
    ,.rlast(merge2_split102_rlast)
    ,.rready(merge2_split102_rready)
    ,.rresp(merge2_split102_rresp[1:0])
    ,.rvalid(merge2_split102_rvalid)
    ,.wdata(merge2_split102_wdata[(DWID - 1):0])
    ,.wlast(merge2_split102_wlast)
    ,.wready(merge2_split102_wready)
    ,.wstrb(merge2_split102_wstrb[(WSTRB - 1):0])
    ,.wvalid(merge2_split102_wvalid)

    ,.a_araddr(split102_merge201_araddr[31:0])
    ,.a_arburst(split102_merge201_arburst[1:0])
    ,.a_arextras(split102_merge201_arextras[(EXTRAS - 1):0])
    ,.a_arid(split102_merge201_arid[(IDWID - 1):0])
    ,.a_arlen(split102_merge201_arlen[7:0])
    ,.a_arready(split102_merge201_arready)
    ,.a_arvalid(split102_merge201_arvalid)
    ,.a_awaddr(split102_merge201_awaddr[31:0])
    ,.a_awburst(split102_merge201_awburst[1:0])
    ,.a_awextras(split102_merge201_awextras[(EXTRAS - 1):0])
    ,.a_awid(split102_merge201_awid[(IDWID - 1):0])
    ,.a_awlen(split102_merge201_awlen[7:0])
    ,.a_awready(split102_merge201_awready)
    ,.a_awvalid(split102_merge201_awvalid)
    ,.a_bid(split102_merge201_bid[(IDWID - 1):0])
    ,.a_bready(split102_merge201_bready)
    ,.a_bresp(split102_merge201_bresp[1:0])
    ,.a_bvalid(split102_merge201_bvalid)
    ,.a_rdata(split102_merge201_rdata[(DWID - 1):0])
    ,.a_rid(split102_merge201_rid[(IDWID - 1):0])
    ,.a_rlast(split102_merge201_rlast)
    ,.a_rready(split102_merge201_rready)
    ,.a_rresp(split102_merge201_rresp[1:0])
    ,.a_rvalid(split102_merge201_rvalid)
    ,.a_wdata(split102_merge201_wdata[(DWID - 1):0])
    ,.a_wlast(split102_merge201_wlast)
    ,.a_wready(split102_merge201_wready)
    ,.a_wstrb(split102_merge201_wstrb[(WSTRB - 1):0])
    ,.a_wvalid(split102_merge201_wvalid)
    ,.b_araddr(split102_merge200_araddr[31:0])
    ,.b_arburst(split102_merge200_arburst[1:0])
    ,.b_arextras(split102_merge200_arextras[(EXTRAS - 1):0])
    ,.b_arid(split102_merge200_arid[(IDWID - 1):0])
    ,.b_arlen(split102_merge200_arlen[7:0])
    ,.b_arready(split102_merge200_arready)
    ,.b_arvalid(split102_merge200_arvalid)
    ,.b_awaddr(split102_merge200_awaddr[31:0])
    ,.b_awburst(split102_merge200_awburst[1:0])
    ,.b_awextras(split102_merge200_awextras[(EXTRAS - 1):0])
    ,.b_awid(split102_merge200_awid[(IDWID - 1):0])
    ,.b_awlen(split102_merge200_awlen[7:0])
    ,.b_awready(split102_merge200_awready)
    ,.b_awvalid(split102_merge200_awvalid)
    ,.b_bid(split102_merge200_bid[(IDWID - 1):0])
    ,.b_bready(split102_merge200_bready)
    ,.b_bresp(split102_merge200_bresp[1:0])
    ,.b_bvalid(split102_merge200_bvalid)
    ,.b_rdata(split102_merge200_rdata[(DWID - 1):0])
    ,.b_rid(split102_merge200_rid[(IDWID - 1):0])
    ,.b_rlast(split102_merge200_rlast)
    ,.b_rready(split102_merge200_rready)
    ,.b_rresp(split102_merge200_rresp[1:0])
    ,.b_rvalid(split102_merge200_rvalid)
    ,.b_wdata(split102_merge200_wdata[(DWID - 1):0])
    ,.b_wlast(split102_merge200_wlast)
    ,.b_wready(split102_merge200_wready)
    ,.b_wstrb(split102_merge200_wstrb[(WSTRB - 1):0])
    ,.b_wvalid(split102_merge200_wvalid)
    ,.c_araddr(split102_merge207_araddr[31:0])
    ,.c_arburst(split102_merge207_arburst[1:0])
    ,.c_arextras(split102_merge207_arextras[(EXTRAS - 1):0])
    ,.c_arid(split102_merge207_arid[(IDWID - 1):0])
    ,.c_arlen(split102_merge207_arlen[7:0])
    ,.c_arready(split102_merge207_arready)
    ,.c_arvalid(split102_merge207_arvalid)
    ,.c_awaddr(split102_merge207_awaddr[31:0])
    ,.c_awburst(split102_merge207_awburst[1:0])
    ,.c_awextras(split102_merge207_awextras[(EXTRAS - 1):0])
    ,.c_awid(split102_merge207_awid[(IDWID - 1):0])
    ,.c_awlen(split102_merge207_awlen[7:0])
    ,.c_awready(split102_merge207_awready)
    ,.c_awvalid(split102_merge207_awvalid)
    ,.c_bid(split102_merge207_bid[(IDWID - 1):0])
    ,.c_bready(split102_merge207_bready)
    ,.c_bresp(split102_merge207_bresp[1:0])
    ,.c_bvalid(split102_merge207_bvalid)
    ,.c_rdata(split102_merge207_rdata[(DWID - 1):0])
    ,.c_rid(split102_merge207_rid[(IDWID - 1):0])
    ,.c_rlast(split102_merge207_rlast)
    ,.c_rready(split102_merge207_rready)
    ,.c_rresp(split102_merge207_rresp[1:0])
    ,.c_rvalid(split102_merge207_rvalid)
    ,.c_wdata(split102_merge207_wdata[(DWID - 1):0])
    ,.c_wlast(split102_merge207_wlast)
    ,.c_wready(split102_merge207_wready)
    ,.c_wstrb(split102_merge207_wstrb[(WSTRB - 1):0])
    ,.c_wvalid(split102_merge207_wvalid)
    ,.d_araddr(split102_merge205_araddr[31:0])
    ,.d_arburst(split102_merge205_arburst[1:0])
    ,.d_arextras(split102_merge205_arextras[(EXTRAS - 1):0])
    ,.d_arid(split102_merge205_arid[(IDWID - 1):0])
    ,.d_arlen(split102_merge205_arlen[7:0])
    ,.d_arready(split102_merge205_arready)
    ,.d_arvalid(split102_merge205_arvalid)
    ,.d_awaddr(split102_merge205_awaddr[31:0])
    ,.d_awburst(split102_merge205_awburst[1:0])
    ,.d_awextras(split102_merge205_awextras[(EXTRAS - 1):0])
    ,.d_awid(split102_merge205_awid[(IDWID - 1):0])
    ,.d_awlen(split102_merge205_awlen[7:0])
    ,.d_awready(split102_merge205_awready)
    ,.d_awvalid(split102_merge205_awvalid)
    ,.d_bid(split102_merge205_bid[(IDWID - 1):0])
    ,.d_bready(split102_merge205_bready)
    ,.d_bresp(split102_merge205_bresp[1:0])
    ,.d_bvalid(split102_merge205_bvalid)
    ,.d_rdata(split102_merge205_rdata[(DWID - 1):0])
    ,.d_rid(split102_merge205_rid[(IDWID - 1):0])
    ,.d_rlast(split102_merge205_rlast)
    ,.d_rready(split102_merge205_rready)
    ,.d_rresp(split102_merge205_rresp[1:0])
    ,.d_rvalid(split102_merge205_rvalid)
    ,.d_wdata(split102_merge205_wdata[(DWID - 1):0])
    ,.d_wlast(split102_merge205_wlast)
    ,.d_wready(split102_merge205_wready)
    ,.d_wstrb(split102_merge205_wstrb[(WSTRB - 1):0])
    ,.d_wvalid(split102_merge205_wvalid)

);

wire [IDWID-1:0] split103_merge200_arid ;
wire [31:0] split103_merge200_araddr ;
wire [7:0] split103_merge200_arlen ;
wire [EXTRAS-1:0] split103_merge200_arextras ;
wire [1:0] split103_merge200_arburst ;
wire split103_merge200_arvalid ;
wire split103_merge200_arready ;
wire [IDWID-1:0] split103_merge200_rid ;
wire [DWID-1:0] split103_merge200_rdata ;
wire [1:0] split103_merge200_rresp ;
wire split103_merge200_rlast ;
wire split103_merge200_rvalid ;
wire split103_merge200_rready ;

wire [IDWID-1:0] split103_merge200_awid ;
wire [31:0] split103_merge200_awaddr ;
wire [7:0] split103_merge200_awlen ;
wire [EXTRAS-1:0] split103_merge200_awextras ;
wire [1:0] split103_merge200_awburst ;
wire split103_merge200_awvalid ;
wire split103_merge200_awready ;
wire [DWID-1:0] split103_merge200_wdata ;
wire [WSTRB-1:0] split103_merge200_wstrb ;
wire split103_merge200_wlast ;
wire split103_merge200_wvalid ;
wire split103_merge200_wready ;
wire [IDWID-1:0] split103_merge200_bid ;
wire [1:0] split103_merge200_bresp ;
wire split103_merge200_bvalid ;
wire split103_merge200_bready ;


wire [IDWID-1:0] split103_merge207_arid ;
wire [31:0] split103_merge207_araddr ;
wire [7:0] split103_merge207_arlen ;
wire [EXTRAS-1:0] split103_merge207_arextras ;
wire [1:0] split103_merge207_arburst ;
wire split103_merge207_arvalid ;
wire split103_merge207_arready ;
wire [IDWID-1:0] split103_merge207_rid ;
wire [DWID-1:0] split103_merge207_rdata ;
wire [1:0] split103_merge207_rresp ;
wire split103_merge207_rlast ;
wire split103_merge207_rvalid ;
wire split103_merge207_rready ;

wire [IDWID-1:0] split103_merge207_awid ;
wire [31:0] split103_merge207_awaddr ;
wire [7:0] split103_merge207_awlen ;
wire [EXTRAS-1:0] split103_merge207_awextras ;
wire [1:0] split103_merge207_awburst ;
wire split103_merge207_awvalid ;
wire split103_merge207_awready ;
wire [DWID-1:0] split103_merge207_wdata ;
wire [WSTRB-1:0] split103_merge207_wstrb ;
wire split103_merge207_wlast ;
wire split103_merge207_wvalid ;
wire split103_merge207_wready ;
wire [IDWID-1:0] split103_merge207_bid ;
wire [1:0] split103_merge207_bresp ;
wire split103_merge207_bvalid ;
wire split103_merge207_bready ;


wire [IDWID-1:0] split103_merge206_arid ;
wire [31:0] split103_merge206_araddr ;
wire [7:0] split103_merge206_arlen ;
wire [EXTRAS-1:0] split103_merge206_arextras ;
wire [1:0] split103_merge206_arburst ;
wire split103_merge206_arvalid ;
wire split103_merge206_arready ;
wire [IDWID-1:0] split103_merge206_rid ;
wire [DWID-1:0] split103_merge206_rdata ;
wire [1:0] split103_merge206_rresp ;
wire split103_merge206_rlast ;
wire split103_merge206_rvalid ;
wire split103_merge206_rready ;

wire [IDWID-1:0] split103_merge206_awid ;
wire [31:0] split103_merge206_awaddr ;
wire [7:0] split103_merge206_awlen ;
wire [EXTRAS-1:0] split103_merge206_awextras ;
wire [1:0] split103_merge206_awburst ;
wire split103_merge206_awvalid ;
wire split103_merge206_awready ;
wire [DWID-1:0] split103_merge206_wdata ;
wire [WSTRB-1:0] split103_merge206_wstrb ;
wire split103_merge206_wlast ;
wire split103_merge206_wvalid ;
wire split103_merge206_wready ;
wire [IDWID-1:0] split103_merge206_bid ;
wire [1:0] split103_merge206_bresp ;
wire split103_merge206_bvalid ;
wire split103_merge206_bready ;


wire [IDWID-1:0] split103_merge203_arid ;
wire [31:0] split103_merge203_araddr ;
wire [7:0] split103_merge203_arlen ;
wire [EXTRAS-1:0] split103_merge203_arextras ;
wire [1:0] split103_merge203_arburst ;
wire split103_merge203_arvalid ;
wire split103_merge203_arready ;
wire [IDWID-1:0] split103_merge203_rid ;
wire [DWID-1:0] split103_merge203_rdata ;
wire [1:0] split103_merge203_rresp ;
wire split103_merge203_rlast ;
wire split103_merge203_rvalid ;
wire split103_merge203_rready ;

wire [IDWID-1:0] split103_merge203_awid ;
wire [31:0] split103_merge203_awaddr ;
wire [7:0] split103_merge203_awlen ;
wire [EXTRAS-1:0] split103_merge203_awextras ;
wire [1:0] split103_merge203_awburst ;
wire split103_merge203_awvalid ;
wire split103_merge203_awready ;
wire [DWID-1:0] split103_merge203_wdata ;
wire [WSTRB-1:0] split103_merge203_wstrb ;
wire split103_merge203_wlast ;
wire split103_merge203_wvalid ;
wire split103_merge203_wready ;
wire [IDWID-1:0] split103_merge203_bid ;
wire [1:0] split103_merge203_bresp ;
wire split103_merge203_bvalid ;
wire split103_merge203_bready ;


axi_4_splitter split103 (
     .clk(clk) ,.rst_n(rst_n)

    ,.araddr(merge3_split103_araddr[31:0])
    ,.arburst(merge3_split103_arburst[1:0])
    ,.arextras(merge3_split103_arextras[(EXTRAS - 1):0])
    ,.arid(merge3_split103_arid[(IDWID - 1):0])
    ,.arlen(merge3_split103_arlen[7:0])
    ,.arready(merge3_split103_arready)
    ,.arvalid(merge3_split103_arvalid)
    ,.awaddr(merge3_split103_awaddr[31:0])
    ,.awburst(merge3_split103_awburst[1:0])
    ,.awextras(merge3_split103_awextras[(EXTRAS - 1):0])
    ,.awid(merge3_split103_awid[3:0])
    ,.awlen(merge3_split103_awlen[7:0])
    ,.awready(merge3_split103_awready)
    ,.awvalid(merge3_split103_awvalid)
    ,.bid(merge3_split103_bid[(IDWID - 1):0])
    ,.bready(merge3_split103_bready)
    ,.bresp(merge3_split103_bresp[1:0])
    ,.bvalid(merge3_split103_bvalid)
    ,.rdata(merge3_split103_rdata[(DWID - 1):0])
    ,.rid(merge3_split103_rid[(IDWID - 1):0])
    ,.rlast(merge3_split103_rlast)
    ,.rready(merge3_split103_rready)
    ,.rresp(merge3_split103_rresp[1:0])
    ,.rvalid(merge3_split103_rvalid)
    ,.wdata(merge3_split103_wdata[(DWID - 1):0])
    ,.wlast(merge3_split103_wlast)
    ,.wready(merge3_split103_wready)
    ,.wstrb(merge3_split103_wstrb[(WSTRB - 1):0])
    ,.wvalid(merge3_split103_wvalid)

    ,.a_araddr(split103_merge200_araddr[31:0])
    ,.a_arburst(split103_merge200_arburst[1:0])
    ,.a_arextras(split103_merge200_arextras[(EXTRAS - 1):0])
    ,.a_arid(split103_merge200_arid[(IDWID - 1):0])
    ,.a_arlen(split103_merge200_arlen[7:0])
    ,.a_arready(split103_merge200_arready)
    ,.a_arvalid(split103_merge200_arvalid)
    ,.a_awaddr(split103_merge200_awaddr[31:0])
    ,.a_awburst(split103_merge200_awburst[1:0])
    ,.a_awextras(split103_merge200_awextras[(EXTRAS - 1):0])
    ,.a_awid(split103_merge200_awid[(IDWID - 1):0])
    ,.a_awlen(split103_merge200_awlen[7:0])
    ,.a_awready(split103_merge200_awready)
    ,.a_awvalid(split103_merge200_awvalid)
    ,.a_bid(split103_merge200_bid[(IDWID - 1):0])
    ,.a_bready(split103_merge200_bready)
    ,.a_bresp(split103_merge200_bresp[1:0])
    ,.a_bvalid(split103_merge200_bvalid)
    ,.a_rdata(split103_merge200_rdata[(DWID - 1):0])
    ,.a_rid(split103_merge200_rid[(IDWID - 1):0])
    ,.a_rlast(split103_merge200_rlast)
    ,.a_rready(split103_merge200_rready)
    ,.a_rresp(split103_merge200_rresp[1:0])
    ,.a_rvalid(split103_merge200_rvalid)
    ,.a_wdata(split103_merge200_wdata[(DWID - 1):0])
    ,.a_wlast(split103_merge200_wlast)
    ,.a_wready(split103_merge200_wready)
    ,.a_wstrb(split103_merge200_wstrb[(WSTRB - 1):0])
    ,.a_wvalid(split103_merge200_wvalid)
    ,.b_araddr(split103_merge207_araddr[31:0])
    ,.b_arburst(split103_merge207_arburst[1:0])
    ,.b_arextras(split103_merge207_arextras[(EXTRAS - 1):0])
    ,.b_arid(split103_merge207_arid[(IDWID - 1):0])
    ,.b_arlen(split103_merge207_arlen[7:0])
    ,.b_arready(split103_merge207_arready)
    ,.b_arvalid(split103_merge207_arvalid)
    ,.b_awaddr(split103_merge207_awaddr[31:0])
    ,.b_awburst(split103_merge207_awburst[1:0])
    ,.b_awextras(split103_merge207_awextras[(EXTRAS - 1):0])
    ,.b_awid(split103_merge207_awid[(IDWID - 1):0])
    ,.b_awlen(split103_merge207_awlen[7:0])
    ,.b_awready(split103_merge207_awready)
    ,.b_awvalid(split103_merge207_awvalid)
    ,.b_bid(split103_merge207_bid[(IDWID - 1):0])
    ,.b_bready(split103_merge207_bready)
    ,.b_bresp(split103_merge207_bresp[1:0])
    ,.b_bvalid(split103_merge207_bvalid)
    ,.b_rdata(split103_merge207_rdata[(DWID - 1):0])
    ,.b_rid(split103_merge207_rid[(IDWID - 1):0])
    ,.b_rlast(split103_merge207_rlast)
    ,.b_rready(split103_merge207_rready)
    ,.b_rresp(split103_merge207_rresp[1:0])
    ,.b_rvalid(split103_merge207_rvalid)
    ,.b_wdata(split103_merge207_wdata[(DWID - 1):0])
    ,.b_wlast(split103_merge207_wlast)
    ,.b_wready(split103_merge207_wready)
    ,.b_wstrb(split103_merge207_wstrb[(WSTRB - 1):0])
    ,.b_wvalid(split103_merge207_wvalid)
    ,.c_araddr(split103_merge206_araddr[31:0])
    ,.c_arburst(split103_merge206_arburst[1:0])
    ,.c_arextras(split103_merge206_arextras[(EXTRAS - 1):0])
    ,.c_arid(split103_merge206_arid[(IDWID - 1):0])
    ,.c_arlen(split103_merge206_arlen[7:0])
    ,.c_arready(split103_merge206_arready)
    ,.c_arvalid(split103_merge206_arvalid)
    ,.c_awaddr(split103_merge206_awaddr[31:0])
    ,.c_awburst(split103_merge206_awburst[1:0])
    ,.c_awextras(split103_merge206_awextras[(EXTRAS - 1):0])
    ,.c_awid(split103_merge206_awid[(IDWID - 1):0])
    ,.c_awlen(split103_merge206_awlen[7:0])
    ,.c_awready(split103_merge206_awready)
    ,.c_awvalid(split103_merge206_awvalid)
    ,.c_bid(split103_merge206_bid[(IDWID - 1):0])
    ,.c_bready(split103_merge206_bready)
    ,.c_bresp(split103_merge206_bresp[1:0])
    ,.c_bvalid(split103_merge206_bvalid)
    ,.c_rdata(split103_merge206_rdata[(DWID - 1):0])
    ,.c_rid(split103_merge206_rid[(IDWID - 1):0])
    ,.c_rlast(split103_merge206_rlast)
    ,.c_rready(split103_merge206_rready)
    ,.c_rresp(split103_merge206_rresp[1:0])
    ,.c_rvalid(split103_merge206_rvalid)
    ,.c_wdata(split103_merge206_wdata[(DWID - 1):0])
    ,.c_wlast(split103_merge206_wlast)
    ,.c_wready(split103_merge206_wready)
    ,.c_wstrb(split103_merge206_wstrb[(WSTRB - 1):0])
    ,.c_wvalid(split103_merge206_wvalid)
    ,.d_araddr(split103_merge203_araddr[31:0])
    ,.d_arburst(split103_merge203_arburst[1:0])
    ,.d_arextras(split103_merge203_arextras[(EXTRAS - 1):0])
    ,.d_arid(split103_merge203_arid[(IDWID - 1):0])
    ,.d_arlen(split103_merge203_arlen[7:0])
    ,.d_arready(split103_merge203_arready)
    ,.d_arvalid(split103_merge203_arvalid)
    ,.d_awaddr(split103_merge203_awaddr[31:0])
    ,.d_awburst(split103_merge203_awburst[1:0])
    ,.d_awextras(split103_merge203_awextras[(EXTRAS - 1):0])
    ,.d_awid(split103_merge203_awid[(IDWID - 1):0])
    ,.d_awlen(split103_merge203_awlen[7:0])
    ,.d_awready(split103_merge203_awready)
    ,.d_awvalid(split103_merge203_awvalid)
    ,.d_bid(split103_merge203_bid[(IDWID - 1):0])
    ,.d_bready(split103_merge203_bready)
    ,.d_bresp(split103_merge203_bresp[1:0])
    ,.d_bvalid(split103_merge203_bvalid)
    ,.d_rdata(split103_merge203_rdata[(DWID - 1):0])
    ,.d_rid(split103_merge203_rid[(IDWID - 1):0])
    ,.d_rlast(split103_merge203_rlast)
    ,.d_rready(split103_merge203_rready)
    ,.d_rresp(split103_merge203_rresp[1:0])
    ,.d_rvalid(split103_merge203_rvalid)
    ,.d_wdata(split103_merge203_wdata[(DWID - 1):0])
    ,.d_wlast(split103_merge203_wlast)
    ,.d_wready(split103_merge203_wready)
    ,.d_wstrb(split103_merge203_wstrb[(WSTRB - 1):0])
    ,.d_wvalid(split103_merge203_wvalid)

);

wire [IDWID-1:0] split104_merge209_arid ;
wire [31:0] split104_merge209_araddr ;
wire [7:0] split104_merge209_arlen ;
wire [EXTRAS-1:0] split104_merge209_arextras ;
wire [1:0] split104_merge209_arburst ;
wire split104_merge209_arvalid ;
wire split104_merge209_arready ;
wire [IDWID-1:0] split104_merge209_rid ;
wire [DWID-1:0] split104_merge209_rdata ;
wire [1:0] split104_merge209_rresp ;
wire split104_merge209_rlast ;
wire split104_merge209_rvalid ;
wire split104_merge209_rready ;

wire [IDWID-1:0] split104_merge209_awid ;
wire [31:0] split104_merge209_awaddr ;
wire [7:0] split104_merge209_awlen ;
wire [EXTRAS-1:0] split104_merge209_awextras ;
wire [1:0] split104_merge209_awburst ;
wire split104_merge209_awvalid ;
wire split104_merge209_awready ;
wire [DWID-1:0] split104_merge209_wdata ;
wire [WSTRB-1:0] split104_merge209_wstrb ;
wire split104_merge209_wlast ;
wire split104_merge209_wvalid ;
wire split104_merge209_wready ;
wire [IDWID-1:0] split104_merge209_bid ;
wire [1:0] split104_merge209_bresp ;
wire split104_merge209_bvalid ;
wire split104_merge209_bready ;


wire [IDWID-1:0] split104_merge206_arid ;
wire [31:0] split104_merge206_araddr ;
wire [7:0] split104_merge206_arlen ;
wire [EXTRAS-1:0] split104_merge206_arextras ;
wire [1:0] split104_merge206_arburst ;
wire split104_merge206_arvalid ;
wire split104_merge206_arready ;
wire [IDWID-1:0] split104_merge206_rid ;
wire [DWID-1:0] split104_merge206_rdata ;
wire [1:0] split104_merge206_rresp ;
wire split104_merge206_rlast ;
wire split104_merge206_rvalid ;
wire split104_merge206_rready ;

wire [IDWID-1:0] split104_merge206_awid ;
wire [31:0] split104_merge206_awaddr ;
wire [7:0] split104_merge206_awlen ;
wire [EXTRAS-1:0] split104_merge206_awextras ;
wire [1:0] split104_merge206_awburst ;
wire split104_merge206_awvalid ;
wire split104_merge206_awready ;
wire [DWID-1:0] split104_merge206_wdata ;
wire [WSTRB-1:0] split104_merge206_wstrb ;
wire split104_merge206_wlast ;
wire split104_merge206_wvalid ;
wire split104_merge206_wready ;
wire [IDWID-1:0] split104_merge206_bid ;
wire [1:0] split104_merge206_bresp ;
wire split104_merge206_bvalid ;
wire split104_merge206_bready ;


wire [IDWID-1:0] split104_merge213_arid ;
wire [31:0] split104_merge213_araddr ;
wire [7:0] split104_merge213_arlen ;
wire [EXTRAS-1:0] split104_merge213_arextras ;
wire [1:0] split104_merge213_arburst ;
wire split104_merge213_arvalid ;
wire split104_merge213_arready ;
wire [IDWID-1:0] split104_merge213_rid ;
wire [DWID-1:0] split104_merge213_rdata ;
wire [1:0] split104_merge213_rresp ;
wire split104_merge213_rlast ;
wire split104_merge213_rvalid ;
wire split104_merge213_rready ;

wire [IDWID-1:0] split104_merge213_awid ;
wire [31:0] split104_merge213_awaddr ;
wire [7:0] split104_merge213_awlen ;
wire [EXTRAS-1:0] split104_merge213_awextras ;
wire [1:0] split104_merge213_awburst ;
wire split104_merge213_awvalid ;
wire split104_merge213_awready ;
wire [DWID-1:0] split104_merge213_wdata ;
wire [WSTRB-1:0] split104_merge213_wstrb ;
wire split104_merge213_wlast ;
wire split104_merge213_wvalid ;
wire split104_merge213_wready ;
wire [IDWID-1:0] split104_merge213_bid ;
wire [1:0] split104_merge213_bresp ;
wire split104_merge213_bvalid ;
wire split104_merge213_bready ;


wire [IDWID-1:0] split104_merge214_arid ;
wire [31:0] split104_merge214_araddr ;
wire [7:0] split104_merge214_arlen ;
wire [EXTRAS-1:0] split104_merge214_arextras ;
wire [1:0] split104_merge214_arburst ;
wire split104_merge214_arvalid ;
wire split104_merge214_arready ;
wire [IDWID-1:0] split104_merge214_rid ;
wire [DWID-1:0] split104_merge214_rdata ;
wire [1:0] split104_merge214_rresp ;
wire split104_merge214_rlast ;
wire split104_merge214_rvalid ;
wire split104_merge214_rready ;

wire [IDWID-1:0] split104_merge214_awid ;
wire [31:0] split104_merge214_awaddr ;
wire [7:0] split104_merge214_awlen ;
wire [EXTRAS-1:0] split104_merge214_awextras ;
wire [1:0] split104_merge214_awburst ;
wire split104_merge214_awvalid ;
wire split104_merge214_awready ;
wire [DWID-1:0] split104_merge214_wdata ;
wire [WSTRB-1:0] split104_merge214_wstrb ;
wire split104_merge214_wlast ;
wire split104_merge214_wvalid ;
wire split104_merge214_wready ;
wire [IDWID-1:0] split104_merge214_bid ;
wire [1:0] split104_merge214_bresp ;
wire split104_merge214_bvalid ;
wire split104_merge214_bready ;


axi_4_splitter split104 (
     .clk(clk) ,.rst_n(rst_n)

    ,.araddr(merge4_split104_araddr[31:0])
    ,.arburst(merge4_split104_arburst[1:0])
    ,.arextras(merge4_split104_arextras[(EXTRAS - 1):0])
    ,.arid(merge4_split104_arid[(IDWID - 1):0])
    ,.arlen(merge4_split104_arlen[7:0])
    ,.arready(merge4_split104_arready)
    ,.arvalid(merge4_split104_arvalid)
    ,.awaddr(merge4_split104_awaddr[31:0])
    ,.awburst(merge4_split104_awburst[1:0])
    ,.awextras(merge4_split104_awextras[(EXTRAS - 1):0])
    ,.awid(merge4_split104_awid[3:0])
    ,.awlen(merge4_split104_awlen[7:0])
    ,.awready(merge4_split104_awready)
    ,.awvalid(merge4_split104_awvalid)
    ,.bid(merge4_split104_bid[(IDWID - 1):0])
    ,.bready(merge4_split104_bready)
    ,.bresp(merge4_split104_bresp[1:0])
    ,.bvalid(merge4_split104_bvalid)
    ,.rdata(merge4_split104_rdata[(DWID - 1):0])
    ,.rid(merge4_split104_rid[(IDWID - 1):0])
    ,.rlast(merge4_split104_rlast)
    ,.rready(merge4_split104_rready)
    ,.rresp(merge4_split104_rresp[1:0])
    ,.rvalid(merge4_split104_rvalid)
    ,.wdata(merge4_split104_wdata[(DWID - 1):0])
    ,.wlast(merge4_split104_wlast)
    ,.wready(merge4_split104_wready)
    ,.wstrb(merge4_split104_wstrb[(WSTRB - 1):0])
    ,.wvalid(merge4_split104_wvalid)

    ,.a_araddr(split104_merge209_araddr[31:0])
    ,.a_arburst(split104_merge209_arburst[1:0])
    ,.a_arextras(split104_merge209_arextras[(EXTRAS - 1):0])
    ,.a_arid(split104_merge209_arid[(IDWID - 1):0])
    ,.a_arlen(split104_merge209_arlen[7:0])
    ,.a_arready(split104_merge209_arready)
    ,.a_arvalid(split104_merge209_arvalid)
    ,.a_awaddr(split104_merge209_awaddr[31:0])
    ,.a_awburst(split104_merge209_awburst[1:0])
    ,.a_awextras(split104_merge209_awextras[(EXTRAS - 1):0])
    ,.a_awid(split104_merge209_awid[(IDWID - 1):0])
    ,.a_awlen(split104_merge209_awlen[7:0])
    ,.a_awready(split104_merge209_awready)
    ,.a_awvalid(split104_merge209_awvalid)
    ,.a_bid(split104_merge209_bid[(IDWID - 1):0])
    ,.a_bready(split104_merge209_bready)
    ,.a_bresp(split104_merge209_bresp[1:0])
    ,.a_bvalid(split104_merge209_bvalid)
    ,.a_rdata(split104_merge209_rdata[(DWID - 1):0])
    ,.a_rid(split104_merge209_rid[(IDWID - 1):0])
    ,.a_rlast(split104_merge209_rlast)
    ,.a_rready(split104_merge209_rready)
    ,.a_rresp(split104_merge209_rresp[1:0])
    ,.a_rvalid(split104_merge209_rvalid)
    ,.a_wdata(split104_merge209_wdata[(DWID - 1):0])
    ,.a_wlast(split104_merge209_wlast)
    ,.a_wready(split104_merge209_wready)
    ,.a_wstrb(split104_merge209_wstrb[(WSTRB - 1):0])
    ,.a_wvalid(split104_merge209_wvalid)
    ,.b_araddr(split104_merge206_araddr[31:0])
    ,.b_arburst(split104_merge206_arburst[1:0])
    ,.b_arextras(split104_merge206_arextras[(EXTRAS - 1):0])
    ,.b_arid(split104_merge206_arid[(IDWID - 1):0])
    ,.b_arlen(split104_merge206_arlen[7:0])
    ,.b_arready(split104_merge206_arready)
    ,.b_arvalid(split104_merge206_arvalid)
    ,.b_awaddr(split104_merge206_awaddr[31:0])
    ,.b_awburst(split104_merge206_awburst[1:0])
    ,.b_awextras(split104_merge206_awextras[(EXTRAS - 1):0])
    ,.b_awid(split104_merge206_awid[(IDWID - 1):0])
    ,.b_awlen(split104_merge206_awlen[7:0])
    ,.b_awready(split104_merge206_awready)
    ,.b_awvalid(split104_merge206_awvalid)
    ,.b_bid(split104_merge206_bid[(IDWID - 1):0])
    ,.b_bready(split104_merge206_bready)
    ,.b_bresp(split104_merge206_bresp[1:0])
    ,.b_bvalid(split104_merge206_bvalid)
    ,.b_rdata(split104_merge206_rdata[(DWID - 1):0])
    ,.b_rid(split104_merge206_rid[(IDWID - 1):0])
    ,.b_rlast(split104_merge206_rlast)
    ,.b_rready(split104_merge206_rready)
    ,.b_rresp(split104_merge206_rresp[1:0])
    ,.b_rvalid(split104_merge206_rvalid)
    ,.b_wdata(split104_merge206_wdata[(DWID - 1):0])
    ,.b_wlast(split104_merge206_wlast)
    ,.b_wready(split104_merge206_wready)
    ,.b_wstrb(split104_merge206_wstrb[(WSTRB - 1):0])
    ,.b_wvalid(split104_merge206_wvalid)
    ,.c_araddr(split104_merge213_araddr[31:0])
    ,.c_arburst(split104_merge213_arburst[1:0])
    ,.c_arextras(split104_merge213_arextras[(EXTRAS - 1):0])
    ,.c_arid(split104_merge213_arid[(IDWID - 1):0])
    ,.c_arlen(split104_merge213_arlen[7:0])
    ,.c_arready(split104_merge213_arready)
    ,.c_arvalid(split104_merge213_arvalid)
    ,.c_awaddr(split104_merge213_awaddr[31:0])
    ,.c_awburst(split104_merge213_awburst[1:0])
    ,.c_awextras(split104_merge213_awextras[(EXTRAS - 1):0])
    ,.c_awid(split104_merge213_awid[(IDWID - 1):0])
    ,.c_awlen(split104_merge213_awlen[7:0])
    ,.c_awready(split104_merge213_awready)
    ,.c_awvalid(split104_merge213_awvalid)
    ,.c_bid(split104_merge213_bid[(IDWID - 1):0])
    ,.c_bready(split104_merge213_bready)
    ,.c_bresp(split104_merge213_bresp[1:0])
    ,.c_bvalid(split104_merge213_bvalid)
    ,.c_rdata(split104_merge213_rdata[(DWID - 1):0])
    ,.c_rid(split104_merge213_rid[(IDWID - 1):0])
    ,.c_rlast(split104_merge213_rlast)
    ,.c_rready(split104_merge213_rready)
    ,.c_rresp(split104_merge213_rresp[1:0])
    ,.c_rvalid(split104_merge213_rvalid)
    ,.c_wdata(split104_merge213_wdata[(DWID - 1):0])
    ,.c_wlast(split104_merge213_wlast)
    ,.c_wready(split104_merge213_wready)
    ,.c_wstrb(split104_merge213_wstrb[(WSTRB - 1):0])
    ,.c_wvalid(split104_merge213_wvalid)
    ,.d_araddr(split104_merge214_araddr[31:0])
    ,.d_arburst(split104_merge214_arburst[1:0])
    ,.d_arextras(split104_merge214_arextras[(EXTRAS - 1):0])
    ,.d_arid(split104_merge214_arid[(IDWID - 1):0])
    ,.d_arlen(split104_merge214_arlen[7:0])
    ,.d_arready(split104_merge214_arready)
    ,.d_arvalid(split104_merge214_arvalid)
    ,.d_awaddr(split104_merge214_awaddr[31:0])
    ,.d_awburst(split104_merge214_awburst[1:0])
    ,.d_awextras(split104_merge214_awextras[(EXTRAS - 1):0])
    ,.d_awid(split104_merge214_awid[(IDWID - 1):0])
    ,.d_awlen(split104_merge214_awlen[7:0])
    ,.d_awready(split104_merge214_awready)
    ,.d_awvalid(split104_merge214_awvalid)
    ,.d_bid(split104_merge214_bid[(IDWID - 1):0])
    ,.d_bready(split104_merge214_bready)
    ,.d_bresp(split104_merge214_bresp[1:0])
    ,.d_bvalid(split104_merge214_bvalid)
    ,.d_rdata(split104_merge214_rdata[(DWID - 1):0])
    ,.d_rid(split104_merge214_rid[(IDWID - 1):0])
    ,.d_rlast(split104_merge214_rlast)
    ,.d_rready(split104_merge214_rready)
    ,.d_rresp(split104_merge214_rresp[1:0])
    ,.d_rvalid(split104_merge214_rvalid)
    ,.d_wdata(split104_merge214_wdata[(DWID - 1):0])
    ,.d_wlast(split104_merge214_wlast)
    ,.d_wready(split104_merge214_wready)
    ,.d_wstrb(split104_merge214_wstrb[(WSTRB - 1):0])
    ,.d_wvalid(split104_merge214_wvalid)

);

wire [IDWID-1:0] split105_merge213_arid ;
wire [31:0] split105_merge213_araddr ;
wire [7:0] split105_merge213_arlen ;
wire [EXTRAS-1:0] split105_merge213_arextras ;
wire [1:0] split105_merge213_arburst ;
wire split105_merge213_arvalid ;
wire split105_merge213_arready ;
wire [IDWID-1:0] split105_merge213_rid ;
wire [DWID-1:0] split105_merge213_rdata ;
wire [1:0] split105_merge213_rresp ;
wire split105_merge213_rlast ;
wire split105_merge213_rvalid ;
wire split105_merge213_rready ;

wire [IDWID-1:0] split105_merge213_awid ;
wire [31:0] split105_merge213_awaddr ;
wire [7:0] split105_merge213_awlen ;
wire [EXTRAS-1:0] split105_merge213_awextras ;
wire [1:0] split105_merge213_awburst ;
wire split105_merge213_awvalid ;
wire split105_merge213_awready ;
wire [DWID-1:0] split105_merge213_wdata ;
wire [WSTRB-1:0] split105_merge213_wstrb ;
wire split105_merge213_wlast ;
wire split105_merge213_wvalid ;
wire split105_merge213_wready ;
wire [IDWID-1:0] split105_merge213_bid ;
wire [1:0] split105_merge213_bresp ;
wire split105_merge213_bvalid ;
wire split105_merge213_bready ;


wire [IDWID-1:0] split105_merge204_arid ;
wire [31:0] split105_merge204_araddr ;
wire [7:0] split105_merge204_arlen ;
wire [EXTRAS-1:0] split105_merge204_arextras ;
wire [1:0] split105_merge204_arburst ;
wire split105_merge204_arvalid ;
wire split105_merge204_arready ;
wire [IDWID-1:0] split105_merge204_rid ;
wire [DWID-1:0] split105_merge204_rdata ;
wire [1:0] split105_merge204_rresp ;
wire split105_merge204_rlast ;
wire split105_merge204_rvalid ;
wire split105_merge204_rready ;

wire [IDWID-1:0] split105_merge204_awid ;
wire [31:0] split105_merge204_awaddr ;
wire [7:0] split105_merge204_awlen ;
wire [EXTRAS-1:0] split105_merge204_awextras ;
wire [1:0] split105_merge204_awburst ;
wire split105_merge204_awvalid ;
wire split105_merge204_awready ;
wire [DWID-1:0] split105_merge204_wdata ;
wire [WSTRB-1:0] split105_merge204_wstrb ;
wire split105_merge204_wlast ;
wire split105_merge204_wvalid ;
wire split105_merge204_wready ;
wire [IDWID-1:0] split105_merge204_bid ;
wire [1:0] split105_merge204_bresp ;
wire split105_merge204_bvalid ;
wire split105_merge204_bready ;


wire [IDWID-1:0] split105_merge208_arid ;
wire [31:0] split105_merge208_araddr ;
wire [7:0] split105_merge208_arlen ;
wire [EXTRAS-1:0] split105_merge208_arextras ;
wire [1:0] split105_merge208_arburst ;
wire split105_merge208_arvalid ;
wire split105_merge208_arready ;
wire [IDWID-1:0] split105_merge208_rid ;
wire [DWID-1:0] split105_merge208_rdata ;
wire [1:0] split105_merge208_rresp ;
wire split105_merge208_rlast ;
wire split105_merge208_rvalid ;
wire split105_merge208_rready ;

wire [IDWID-1:0] split105_merge208_awid ;
wire [31:0] split105_merge208_awaddr ;
wire [7:0] split105_merge208_awlen ;
wire [EXTRAS-1:0] split105_merge208_awextras ;
wire [1:0] split105_merge208_awburst ;
wire split105_merge208_awvalid ;
wire split105_merge208_awready ;
wire [DWID-1:0] split105_merge208_wdata ;
wire [WSTRB-1:0] split105_merge208_wstrb ;
wire split105_merge208_wlast ;
wire split105_merge208_wvalid ;
wire split105_merge208_wready ;
wire [IDWID-1:0] split105_merge208_bid ;
wire [1:0] split105_merge208_bresp ;
wire split105_merge208_bvalid ;
wire split105_merge208_bready ;


wire [IDWID-1:0] split105_merge212_arid ;
wire [31:0] split105_merge212_araddr ;
wire [7:0] split105_merge212_arlen ;
wire [EXTRAS-1:0] split105_merge212_arextras ;
wire [1:0] split105_merge212_arburst ;
wire split105_merge212_arvalid ;
wire split105_merge212_arready ;
wire [IDWID-1:0] split105_merge212_rid ;
wire [DWID-1:0] split105_merge212_rdata ;
wire [1:0] split105_merge212_rresp ;
wire split105_merge212_rlast ;
wire split105_merge212_rvalid ;
wire split105_merge212_rready ;

wire [IDWID-1:0] split105_merge212_awid ;
wire [31:0] split105_merge212_awaddr ;
wire [7:0] split105_merge212_awlen ;
wire [EXTRAS-1:0] split105_merge212_awextras ;
wire [1:0] split105_merge212_awburst ;
wire split105_merge212_awvalid ;
wire split105_merge212_awready ;
wire [DWID-1:0] split105_merge212_wdata ;
wire [WSTRB-1:0] split105_merge212_wstrb ;
wire split105_merge212_wlast ;
wire split105_merge212_wvalid ;
wire split105_merge212_wready ;
wire [IDWID-1:0] split105_merge212_bid ;
wire [1:0] split105_merge212_bresp ;
wire split105_merge212_bvalid ;
wire split105_merge212_bready ;


axi_4_splitter split105 (
     .clk(clk) ,.rst_n(rst_n)

    ,.araddr(merge5_split105_araddr[31:0])
    ,.arburst(merge5_split105_arburst[1:0])
    ,.arextras(merge5_split105_arextras[(EXTRAS - 1):0])
    ,.arid(merge5_split105_arid[(IDWID - 1):0])
    ,.arlen(merge5_split105_arlen[7:0])
    ,.arready(merge5_split105_arready)
    ,.arvalid(merge5_split105_arvalid)
    ,.awaddr(merge5_split105_awaddr[31:0])
    ,.awburst(merge5_split105_awburst[1:0])
    ,.awextras(merge5_split105_awextras[(EXTRAS - 1):0])
    ,.awid(merge5_split105_awid[3:0])
    ,.awlen(merge5_split105_awlen[7:0])
    ,.awready(merge5_split105_awready)
    ,.awvalid(merge5_split105_awvalid)
    ,.bid(merge5_split105_bid[(IDWID - 1):0])
    ,.bready(merge5_split105_bready)
    ,.bresp(merge5_split105_bresp[1:0])
    ,.bvalid(merge5_split105_bvalid)
    ,.rdata(merge5_split105_rdata[(DWID - 1):0])
    ,.rid(merge5_split105_rid[(IDWID - 1):0])
    ,.rlast(merge5_split105_rlast)
    ,.rready(merge5_split105_rready)
    ,.rresp(merge5_split105_rresp[1:0])
    ,.rvalid(merge5_split105_rvalid)
    ,.wdata(merge5_split105_wdata[(DWID - 1):0])
    ,.wlast(merge5_split105_wlast)
    ,.wready(merge5_split105_wready)
    ,.wstrb(merge5_split105_wstrb[(WSTRB - 1):0])
    ,.wvalid(merge5_split105_wvalid)

    ,.a_araddr(split105_merge213_araddr[31:0])
    ,.a_arburst(split105_merge213_arburst[1:0])
    ,.a_arextras(split105_merge213_arextras[(EXTRAS - 1):0])
    ,.a_arid(split105_merge213_arid[(IDWID - 1):0])
    ,.a_arlen(split105_merge213_arlen[7:0])
    ,.a_arready(split105_merge213_arready)
    ,.a_arvalid(split105_merge213_arvalid)
    ,.a_awaddr(split105_merge213_awaddr[31:0])
    ,.a_awburst(split105_merge213_awburst[1:0])
    ,.a_awextras(split105_merge213_awextras[(EXTRAS - 1):0])
    ,.a_awid(split105_merge213_awid[(IDWID - 1):0])
    ,.a_awlen(split105_merge213_awlen[7:0])
    ,.a_awready(split105_merge213_awready)
    ,.a_awvalid(split105_merge213_awvalid)
    ,.a_bid(split105_merge213_bid[(IDWID - 1):0])
    ,.a_bready(split105_merge213_bready)
    ,.a_bresp(split105_merge213_bresp[1:0])
    ,.a_bvalid(split105_merge213_bvalid)
    ,.a_rdata(split105_merge213_rdata[(DWID - 1):0])
    ,.a_rid(split105_merge213_rid[(IDWID - 1):0])
    ,.a_rlast(split105_merge213_rlast)
    ,.a_rready(split105_merge213_rready)
    ,.a_rresp(split105_merge213_rresp[1:0])
    ,.a_rvalid(split105_merge213_rvalid)
    ,.a_wdata(split105_merge213_wdata[(DWID - 1):0])
    ,.a_wlast(split105_merge213_wlast)
    ,.a_wready(split105_merge213_wready)
    ,.a_wstrb(split105_merge213_wstrb[(WSTRB - 1):0])
    ,.a_wvalid(split105_merge213_wvalid)
    ,.b_araddr(split105_merge204_araddr[31:0])
    ,.b_arburst(split105_merge204_arburst[1:0])
    ,.b_arextras(split105_merge204_arextras[(EXTRAS - 1):0])
    ,.b_arid(split105_merge204_arid[(IDWID - 1):0])
    ,.b_arlen(split105_merge204_arlen[7:0])
    ,.b_arready(split105_merge204_arready)
    ,.b_arvalid(split105_merge204_arvalid)
    ,.b_awaddr(split105_merge204_awaddr[31:0])
    ,.b_awburst(split105_merge204_awburst[1:0])
    ,.b_awextras(split105_merge204_awextras[(EXTRAS - 1):0])
    ,.b_awid(split105_merge204_awid[(IDWID - 1):0])
    ,.b_awlen(split105_merge204_awlen[7:0])
    ,.b_awready(split105_merge204_awready)
    ,.b_awvalid(split105_merge204_awvalid)
    ,.b_bid(split105_merge204_bid[(IDWID - 1):0])
    ,.b_bready(split105_merge204_bready)
    ,.b_bresp(split105_merge204_bresp[1:0])
    ,.b_bvalid(split105_merge204_bvalid)
    ,.b_rdata(split105_merge204_rdata[(DWID - 1):0])
    ,.b_rid(split105_merge204_rid[(IDWID - 1):0])
    ,.b_rlast(split105_merge204_rlast)
    ,.b_rready(split105_merge204_rready)
    ,.b_rresp(split105_merge204_rresp[1:0])
    ,.b_rvalid(split105_merge204_rvalid)
    ,.b_wdata(split105_merge204_wdata[(DWID - 1):0])
    ,.b_wlast(split105_merge204_wlast)
    ,.b_wready(split105_merge204_wready)
    ,.b_wstrb(split105_merge204_wstrb[(WSTRB - 1):0])
    ,.b_wvalid(split105_merge204_wvalid)
    ,.c_araddr(split105_merge208_araddr[31:0])
    ,.c_arburst(split105_merge208_arburst[1:0])
    ,.c_arextras(split105_merge208_arextras[(EXTRAS - 1):0])
    ,.c_arid(split105_merge208_arid[(IDWID - 1):0])
    ,.c_arlen(split105_merge208_arlen[7:0])
    ,.c_arready(split105_merge208_arready)
    ,.c_arvalid(split105_merge208_arvalid)
    ,.c_awaddr(split105_merge208_awaddr[31:0])
    ,.c_awburst(split105_merge208_awburst[1:0])
    ,.c_awextras(split105_merge208_awextras[(EXTRAS - 1):0])
    ,.c_awid(split105_merge208_awid[(IDWID - 1):0])
    ,.c_awlen(split105_merge208_awlen[7:0])
    ,.c_awready(split105_merge208_awready)
    ,.c_awvalid(split105_merge208_awvalid)
    ,.c_bid(split105_merge208_bid[(IDWID - 1):0])
    ,.c_bready(split105_merge208_bready)
    ,.c_bresp(split105_merge208_bresp[1:0])
    ,.c_bvalid(split105_merge208_bvalid)
    ,.c_rdata(split105_merge208_rdata[(DWID - 1):0])
    ,.c_rid(split105_merge208_rid[(IDWID - 1):0])
    ,.c_rlast(split105_merge208_rlast)
    ,.c_rready(split105_merge208_rready)
    ,.c_rresp(split105_merge208_rresp[1:0])
    ,.c_rvalid(split105_merge208_rvalid)
    ,.c_wdata(split105_merge208_wdata[(DWID - 1):0])
    ,.c_wlast(split105_merge208_wlast)
    ,.c_wready(split105_merge208_wready)
    ,.c_wstrb(split105_merge208_wstrb[(WSTRB - 1):0])
    ,.c_wvalid(split105_merge208_wvalid)
    ,.d_araddr(split105_merge212_araddr[31:0])
    ,.d_arburst(split105_merge212_arburst[1:0])
    ,.d_arextras(split105_merge212_arextras[(EXTRAS - 1):0])
    ,.d_arid(split105_merge212_arid[(IDWID - 1):0])
    ,.d_arlen(split105_merge212_arlen[7:0])
    ,.d_arready(split105_merge212_arready)
    ,.d_arvalid(split105_merge212_arvalid)
    ,.d_awaddr(split105_merge212_awaddr[31:0])
    ,.d_awburst(split105_merge212_awburst[1:0])
    ,.d_awextras(split105_merge212_awextras[(EXTRAS - 1):0])
    ,.d_awid(split105_merge212_awid[(IDWID - 1):0])
    ,.d_awlen(split105_merge212_awlen[7:0])
    ,.d_awready(split105_merge212_awready)
    ,.d_awvalid(split105_merge212_awvalid)
    ,.d_bid(split105_merge212_bid[(IDWID - 1):0])
    ,.d_bready(split105_merge212_bready)
    ,.d_bresp(split105_merge212_bresp[1:0])
    ,.d_bvalid(split105_merge212_bvalid)
    ,.d_rdata(split105_merge212_rdata[(DWID - 1):0])
    ,.d_rid(split105_merge212_rid[(IDWID - 1):0])
    ,.d_rlast(split105_merge212_rlast)
    ,.d_rready(split105_merge212_rready)
    ,.d_rresp(split105_merge212_rresp[1:0])
    ,.d_rvalid(split105_merge212_rvalid)
    ,.d_wdata(split105_merge212_wdata[(DWID - 1):0])
    ,.d_wlast(split105_merge212_wlast)
    ,.d_wready(split105_merge212_wready)
    ,.d_wstrb(split105_merge212_wstrb[(WSTRB - 1):0])
    ,.d_wvalid(split105_merge212_wvalid)

);

wire [IDWID-1:0] split106_merge213_arid ;
wire [31:0] split106_merge213_araddr ;
wire [7:0] split106_merge213_arlen ;
wire [EXTRAS-1:0] split106_merge213_arextras ;
wire [1:0] split106_merge213_arburst ;
wire split106_merge213_arvalid ;
wire split106_merge213_arready ;
wire [IDWID-1:0] split106_merge213_rid ;
wire [DWID-1:0] split106_merge213_rdata ;
wire [1:0] split106_merge213_rresp ;
wire split106_merge213_rlast ;
wire split106_merge213_rvalid ;
wire split106_merge213_rready ;

wire [IDWID-1:0] split106_merge213_awid ;
wire [31:0] split106_merge213_awaddr ;
wire [7:0] split106_merge213_awlen ;
wire [EXTRAS-1:0] split106_merge213_awextras ;
wire [1:0] split106_merge213_awburst ;
wire split106_merge213_awvalid ;
wire split106_merge213_awready ;
wire [DWID-1:0] split106_merge213_wdata ;
wire [WSTRB-1:0] split106_merge213_wstrb ;
wire split106_merge213_wlast ;
wire split106_merge213_wvalid ;
wire split106_merge213_wready ;
wire [IDWID-1:0] split106_merge213_bid ;
wire [1:0] split106_merge213_bresp ;
wire split106_merge213_bvalid ;
wire split106_merge213_bready ;


wire [IDWID-1:0] split106_merge205_arid ;
wire [31:0] split106_merge205_araddr ;
wire [7:0] split106_merge205_arlen ;
wire [EXTRAS-1:0] split106_merge205_arextras ;
wire [1:0] split106_merge205_arburst ;
wire split106_merge205_arvalid ;
wire split106_merge205_arready ;
wire [IDWID-1:0] split106_merge205_rid ;
wire [DWID-1:0] split106_merge205_rdata ;
wire [1:0] split106_merge205_rresp ;
wire split106_merge205_rlast ;
wire split106_merge205_rvalid ;
wire split106_merge205_rready ;

wire [IDWID-1:0] split106_merge205_awid ;
wire [31:0] split106_merge205_awaddr ;
wire [7:0] split106_merge205_awlen ;
wire [EXTRAS-1:0] split106_merge205_awextras ;
wire [1:0] split106_merge205_awburst ;
wire split106_merge205_awvalid ;
wire split106_merge205_awready ;
wire [DWID-1:0] split106_merge205_wdata ;
wire [WSTRB-1:0] split106_merge205_wstrb ;
wire split106_merge205_wlast ;
wire split106_merge205_wvalid ;
wire split106_merge205_wready ;
wire [IDWID-1:0] split106_merge205_bid ;
wire [1:0] split106_merge205_bresp ;
wire split106_merge205_bvalid ;
wire split106_merge205_bready ;


wire [IDWID-1:0] split106_merge211_arid ;
wire [31:0] split106_merge211_araddr ;
wire [7:0] split106_merge211_arlen ;
wire [EXTRAS-1:0] split106_merge211_arextras ;
wire [1:0] split106_merge211_arburst ;
wire split106_merge211_arvalid ;
wire split106_merge211_arready ;
wire [IDWID-1:0] split106_merge211_rid ;
wire [DWID-1:0] split106_merge211_rdata ;
wire [1:0] split106_merge211_rresp ;
wire split106_merge211_rlast ;
wire split106_merge211_rvalid ;
wire split106_merge211_rready ;

wire [IDWID-1:0] split106_merge211_awid ;
wire [31:0] split106_merge211_awaddr ;
wire [7:0] split106_merge211_awlen ;
wire [EXTRAS-1:0] split106_merge211_awextras ;
wire [1:0] split106_merge211_awburst ;
wire split106_merge211_awvalid ;
wire split106_merge211_awready ;
wire [DWID-1:0] split106_merge211_wdata ;
wire [WSTRB-1:0] split106_merge211_wstrb ;
wire split106_merge211_wlast ;
wire split106_merge211_wvalid ;
wire split106_merge211_wready ;
wire [IDWID-1:0] split106_merge211_bid ;
wire [1:0] split106_merge211_bresp ;
wire split106_merge211_bvalid ;
wire split106_merge211_bready ;


wire [IDWID-1:0] split106_merge204_arid ;
wire [31:0] split106_merge204_araddr ;
wire [7:0] split106_merge204_arlen ;
wire [EXTRAS-1:0] split106_merge204_arextras ;
wire [1:0] split106_merge204_arburst ;
wire split106_merge204_arvalid ;
wire split106_merge204_arready ;
wire [IDWID-1:0] split106_merge204_rid ;
wire [DWID-1:0] split106_merge204_rdata ;
wire [1:0] split106_merge204_rresp ;
wire split106_merge204_rlast ;
wire split106_merge204_rvalid ;
wire split106_merge204_rready ;

wire [IDWID-1:0] split106_merge204_awid ;
wire [31:0] split106_merge204_awaddr ;
wire [7:0] split106_merge204_awlen ;
wire [EXTRAS-1:0] split106_merge204_awextras ;
wire [1:0] split106_merge204_awburst ;
wire split106_merge204_awvalid ;
wire split106_merge204_awready ;
wire [DWID-1:0] split106_merge204_wdata ;
wire [WSTRB-1:0] split106_merge204_wstrb ;
wire split106_merge204_wlast ;
wire split106_merge204_wvalid ;
wire split106_merge204_wready ;
wire [IDWID-1:0] split106_merge204_bid ;
wire [1:0] split106_merge204_bresp ;
wire split106_merge204_bvalid ;
wire split106_merge204_bready ;


axi_4_splitter split106 (
     .clk(clk) ,.rst_n(rst_n)

    ,.araddr(merge6_split106_araddr[31:0])
    ,.arburst(merge6_split106_arburst[1:0])
    ,.arextras(merge6_split106_arextras[(EXTRAS - 1):0])
    ,.arid(merge6_split106_arid[(IDWID - 1):0])
    ,.arlen(merge6_split106_arlen[7:0])
    ,.arready(merge6_split106_arready)
    ,.arvalid(merge6_split106_arvalid)
    ,.awaddr(merge6_split106_awaddr[31:0])
    ,.awburst(merge6_split106_awburst[1:0])
    ,.awextras(merge6_split106_awextras[(EXTRAS - 1):0])
    ,.awid(merge6_split106_awid[3:0])
    ,.awlen(merge6_split106_awlen[7:0])
    ,.awready(merge6_split106_awready)
    ,.awvalid(merge6_split106_awvalid)
    ,.bid(merge6_split106_bid[(IDWID - 1):0])
    ,.bready(merge6_split106_bready)
    ,.bresp(merge6_split106_bresp[1:0])
    ,.bvalid(merge6_split106_bvalid)
    ,.rdata(merge6_split106_rdata[(DWID - 1):0])
    ,.rid(merge6_split106_rid[(IDWID - 1):0])
    ,.rlast(merge6_split106_rlast)
    ,.rready(merge6_split106_rready)
    ,.rresp(merge6_split106_rresp[1:0])
    ,.rvalid(merge6_split106_rvalid)
    ,.wdata(merge6_split106_wdata[(DWID - 1):0])
    ,.wlast(merge6_split106_wlast)
    ,.wready(merge6_split106_wready)
    ,.wstrb(merge6_split106_wstrb[(WSTRB - 1):0])
    ,.wvalid(merge6_split106_wvalid)

    ,.a_araddr(split106_merge213_araddr[31:0])
    ,.a_arburst(split106_merge213_arburst[1:0])
    ,.a_arextras(split106_merge213_arextras[(EXTRAS - 1):0])
    ,.a_arid(split106_merge213_arid[(IDWID - 1):0])
    ,.a_arlen(split106_merge213_arlen[7:0])
    ,.a_arready(split106_merge213_arready)
    ,.a_arvalid(split106_merge213_arvalid)
    ,.a_awaddr(split106_merge213_awaddr[31:0])
    ,.a_awburst(split106_merge213_awburst[1:0])
    ,.a_awextras(split106_merge213_awextras[(EXTRAS - 1):0])
    ,.a_awid(split106_merge213_awid[(IDWID - 1):0])
    ,.a_awlen(split106_merge213_awlen[7:0])
    ,.a_awready(split106_merge213_awready)
    ,.a_awvalid(split106_merge213_awvalid)
    ,.a_bid(split106_merge213_bid[(IDWID - 1):0])
    ,.a_bready(split106_merge213_bready)
    ,.a_bresp(split106_merge213_bresp[1:0])
    ,.a_bvalid(split106_merge213_bvalid)
    ,.a_rdata(split106_merge213_rdata[(DWID - 1):0])
    ,.a_rid(split106_merge213_rid[(IDWID - 1):0])
    ,.a_rlast(split106_merge213_rlast)
    ,.a_rready(split106_merge213_rready)
    ,.a_rresp(split106_merge213_rresp[1:0])
    ,.a_rvalid(split106_merge213_rvalid)
    ,.a_wdata(split106_merge213_wdata[(DWID - 1):0])
    ,.a_wlast(split106_merge213_wlast)
    ,.a_wready(split106_merge213_wready)
    ,.a_wstrb(split106_merge213_wstrb[(WSTRB - 1):0])
    ,.a_wvalid(split106_merge213_wvalid)
    ,.b_araddr(split106_merge205_araddr[31:0])
    ,.b_arburst(split106_merge205_arburst[1:0])
    ,.b_arextras(split106_merge205_arextras[(EXTRAS - 1):0])
    ,.b_arid(split106_merge205_arid[(IDWID - 1):0])
    ,.b_arlen(split106_merge205_arlen[7:0])
    ,.b_arready(split106_merge205_arready)
    ,.b_arvalid(split106_merge205_arvalid)
    ,.b_awaddr(split106_merge205_awaddr[31:0])
    ,.b_awburst(split106_merge205_awburst[1:0])
    ,.b_awextras(split106_merge205_awextras[(EXTRAS - 1):0])
    ,.b_awid(split106_merge205_awid[(IDWID - 1):0])
    ,.b_awlen(split106_merge205_awlen[7:0])
    ,.b_awready(split106_merge205_awready)
    ,.b_awvalid(split106_merge205_awvalid)
    ,.b_bid(split106_merge205_bid[(IDWID - 1):0])
    ,.b_bready(split106_merge205_bready)
    ,.b_bresp(split106_merge205_bresp[1:0])
    ,.b_bvalid(split106_merge205_bvalid)
    ,.b_rdata(split106_merge205_rdata[(DWID - 1):0])
    ,.b_rid(split106_merge205_rid[(IDWID - 1):0])
    ,.b_rlast(split106_merge205_rlast)
    ,.b_rready(split106_merge205_rready)
    ,.b_rresp(split106_merge205_rresp[1:0])
    ,.b_rvalid(split106_merge205_rvalid)
    ,.b_wdata(split106_merge205_wdata[(DWID - 1):0])
    ,.b_wlast(split106_merge205_wlast)
    ,.b_wready(split106_merge205_wready)
    ,.b_wstrb(split106_merge205_wstrb[(WSTRB - 1):0])
    ,.b_wvalid(split106_merge205_wvalid)
    ,.c_araddr(split106_merge211_araddr[31:0])
    ,.c_arburst(split106_merge211_arburst[1:0])
    ,.c_arextras(split106_merge211_arextras[(EXTRAS - 1):0])
    ,.c_arid(split106_merge211_arid[(IDWID - 1):0])
    ,.c_arlen(split106_merge211_arlen[7:0])
    ,.c_arready(split106_merge211_arready)
    ,.c_arvalid(split106_merge211_arvalid)
    ,.c_awaddr(split106_merge211_awaddr[31:0])
    ,.c_awburst(split106_merge211_awburst[1:0])
    ,.c_awextras(split106_merge211_awextras[(EXTRAS - 1):0])
    ,.c_awid(split106_merge211_awid[(IDWID - 1):0])
    ,.c_awlen(split106_merge211_awlen[7:0])
    ,.c_awready(split106_merge211_awready)
    ,.c_awvalid(split106_merge211_awvalid)
    ,.c_bid(split106_merge211_bid[(IDWID - 1):0])
    ,.c_bready(split106_merge211_bready)
    ,.c_bresp(split106_merge211_bresp[1:0])
    ,.c_bvalid(split106_merge211_bvalid)
    ,.c_rdata(split106_merge211_rdata[(DWID - 1):0])
    ,.c_rid(split106_merge211_rid[(IDWID - 1):0])
    ,.c_rlast(split106_merge211_rlast)
    ,.c_rready(split106_merge211_rready)
    ,.c_rresp(split106_merge211_rresp[1:0])
    ,.c_rvalid(split106_merge211_rvalid)
    ,.c_wdata(split106_merge211_wdata[(DWID - 1):0])
    ,.c_wlast(split106_merge211_wlast)
    ,.c_wready(split106_merge211_wready)
    ,.c_wstrb(split106_merge211_wstrb[(WSTRB - 1):0])
    ,.c_wvalid(split106_merge211_wvalid)
    ,.d_araddr(split106_merge204_araddr[31:0])
    ,.d_arburst(split106_merge204_arburst[1:0])
    ,.d_arextras(split106_merge204_arextras[(EXTRAS - 1):0])
    ,.d_arid(split106_merge204_arid[(IDWID - 1):0])
    ,.d_arlen(split106_merge204_arlen[7:0])
    ,.d_arready(split106_merge204_arready)
    ,.d_arvalid(split106_merge204_arvalid)
    ,.d_awaddr(split106_merge204_awaddr[31:0])
    ,.d_awburst(split106_merge204_awburst[1:0])
    ,.d_awextras(split106_merge204_awextras[(EXTRAS - 1):0])
    ,.d_awid(split106_merge204_awid[(IDWID - 1):0])
    ,.d_awlen(split106_merge204_awlen[7:0])
    ,.d_awready(split106_merge204_awready)
    ,.d_awvalid(split106_merge204_awvalid)
    ,.d_bid(split106_merge204_bid[(IDWID - 1):0])
    ,.d_bready(split106_merge204_bready)
    ,.d_bresp(split106_merge204_bresp[1:0])
    ,.d_bvalid(split106_merge204_bvalid)
    ,.d_rdata(split106_merge204_rdata[(DWID - 1):0])
    ,.d_rid(split106_merge204_rid[(IDWID - 1):0])
    ,.d_rlast(split106_merge204_rlast)
    ,.d_rready(split106_merge204_rready)
    ,.d_rresp(split106_merge204_rresp[1:0])
    ,.d_rvalid(split106_merge204_rvalid)
    ,.d_wdata(split106_merge204_wdata[(DWID - 1):0])
    ,.d_wlast(split106_merge204_wlast)
    ,.d_wready(split106_merge204_wready)
    ,.d_wstrb(split106_merge204_wstrb[(WSTRB - 1):0])
    ,.d_wvalid(split106_merge204_wvalid)

);

wire [IDWID-1:0] split107_merge210_arid ;
wire [31:0] split107_merge210_araddr ;
wire [7:0] split107_merge210_arlen ;
wire [EXTRAS-1:0] split107_merge210_arextras ;
wire [1:0] split107_merge210_arburst ;
wire split107_merge210_arvalid ;
wire split107_merge210_arready ;
wire [IDWID-1:0] split107_merge210_rid ;
wire [DWID-1:0] split107_merge210_rdata ;
wire [1:0] split107_merge210_rresp ;
wire split107_merge210_rlast ;
wire split107_merge210_rvalid ;
wire split107_merge210_rready ;

wire [IDWID-1:0] split107_merge210_awid ;
wire [31:0] split107_merge210_awaddr ;
wire [7:0] split107_merge210_awlen ;
wire [EXTRAS-1:0] split107_merge210_awextras ;
wire [1:0] split107_merge210_awburst ;
wire split107_merge210_awvalid ;
wire split107_merge210_awready ;
wire [DWID-1:0] split107_merge210_wdata ;
wire [WSTRB-1:0] split107_merge210_wstrb ;
wire split107_merge210_wlast ;
wire split107_merge210_wvalid ;
wire split107_merge210_wready ;
wire [IDWID-1:0] split107_merge210_bid ;
wire [1:0] split107_merge210_bresp ;
wire split107_merge210_bvalid ;
wire split107_merge210_bready ;


wire [IDWID-1:0] split107_merge202_arid ;
wire [31:0] split107_merge202_araddr ;
wire [7:0] split107_merge202_arlen ;
wire [EXTRAS-1:0] split107_merge202_arextras ;
wire [1:0] split107_merge202_arburst ;
wire split107_merge202_arvalid ;
wire split107_merge202_arready ;
wire [IDWID-1:0] split107_merge202_rid ;
wire [DWID-1:0] split107_merge202_rdata ;
wire [1:0] split107_merge202_rresp ;
wire split107_merge202_rlast ;
wire split107_merge202_rvalid ;
wire split107_merge202_rready ;

wire [IDWID-1:0] split107_merge202_awid ;
wire [31:0] split107_merge202_awaddr ;
wire [7:0] split107_merge202_awlen ;
wire [EXTRAS-1:0] split107_merge202_awextras ;
wire [1:0] split107_merge202_awburst ;
wire split107_merge202_awvalid ;
wire split107_merge202_awready ;
wire [DWID-1:0] split107_merge202_wdata ;
wire [WSTRB-1:0] split107_merge202_wstrb ;
wire split107_merge202_wlast ;
wire split107_merge202_wvalid ;
wire split107_merge202_wready ;
wire [IDWID-1:0] split107_merge202_bid ;
wire [1:0] split107_merge202_bresp ;
wire split107_merge202_bvalid ;
wire split107_merge202_bready ;


wire [IDWID-1:0] split107_merge207_arid ;
wire [31:0] split107_merge207_araddr ;
wire [7:0] split107_merge207_arlen ;
wire [EXTRAS-1:0] split107_merge207_arextras ;
wire [1:0] split107_merge207_arburst ;
wire split107_merge207_arvalid ;
wire split107_merge207_arready ;
wire [IDWID-1:0] split107_merge207_rid ;
wire [DWID-1:0] split107_merge207_rdata ;
wire [1:0] split107_merge207_rresp ;
wire split107_merge207_rlast ;
wire split107_merge207_rvalid ;
wire split107_merge207_rready ;

wire [IDWID-1:0] split107_merge207_awid ;
wire [31:0] split107_merge207_awaddr ;
wire [7:0] split107_merge207_awlen ;
wire [EXTRAS-1:0] split107_merge207_awextras ;
wire [1:0] split107_merge207_awburst ;
wire split107_merge207_awvalid ;
wire split107_merge207_awready ;
wire [DWID-1:0] split107_merge207_wdata ;
wire [WSTRB-1:0] split107_merge207_wstrb ;
wire split107_merge207_wlast ;
wire split107_merge207_wvalid ;
wire split107_merge207_wready ;
wire [IDWID-1:0] split107_merge207_bid ;
wire [1:0] split107_merge207_bresp ;
wire split107_merge207_bvalid ;
wire split107_merge207_bready ;


wire [IDWID-1:0] split107_merge211_arid ;
wire [31:0] split107_merge211_araddr ;
wire [7:0] split107_merge211_arlen ;
wire [EXTRAS-1:0] split107_merge211_arextras ;
wire [1:0] split107_merge211_arburst ;
wire split107_merge211_arvalid ;
wire split107_merge211_arready ;
wire [IDWID-1:0] split107_merge211_rid ;
wire [DWID-1:0] split107_merge211_rdata ;
wire [1:0] split107_merge211_rresp ;
wire split107_merge211_rlast ;
wire split107_merge211_rvalid ;
wire split107_merge211_rready ;

wire [IDWID-1:0] split107_merge211_awid ;
wire [31:0] split107_merge211_awaddr ;
wire [7:0] split107_merge211_awlen ;
wire [EXTRAS-1:0] split107_merge211_awextras ;
wire [1:0] split107_merge211_awburst ;
wire split107_merge211_awvalid ;
wire split107_merge211_awready ;
wire [DWID-1:0] split107_merge211_wdata ;
wire [WSTRB-1:0] split107_merge211_wstrb ;
wire split107_merge211_wlast ;
wire split107_merge211_wvalid ;
wire split107_merge211_wready ;
wire [IDWID-1:0] split107_merge211_bid ;
wire [1:0] split107_merge211_bresp ;
wire split107_merge211_bvalid ;
wire split107_merge211_bready ;


axi_4_splitter split107 (
     .clk(clk) ,.rst_n(rst_n)

    ,.araddr(merge7_split107_araddr[31:0])
    ,.arburst(merge7_split107_arburst[1:0])
    ,.arextras(merge7_split107_arextras[(EXTRAS - 1):0])
    ,.arid(merge7_split107_arid[(IDWID - 1):0])
    ,.arlen(merge7_split107_arlen[7:0])
    ,.arready(merge7_split107_arready)
    ,.arvalid(merge7_split107_arvalid)
    ,.awaddr(merge7_split107_awaddr[31:0])
    ,.awburst(merge7_split107_awburst[1:0])
    ,.awextras(merge7_split107_awextras[(EXTRAS - 1):0])
    ,.awid(merge7_split107_awid[3:0])
    ,.awlen(merge7_split107_awlen[7:0])
    ,.awready(merge7_split107_awready)
    ,.awvalid(merge7_split107_awvalid)
    ,.bid(merge7_split107_bid[(IDWID - 1):0])
    ,.bready(merge7_split107_bready)
    ,.bresp(merge7_split107_bresp[1:0])
    ,.bvalid(merge7_split107_bvalid)
    ,.rdata(merge7_split107_rdata[(DWID - 1):0])
    ,.rid(merge7_split107_rid[(IDWID - 1):0])
    ,.rlast(merge7_split107_rlast)
    ,.rready(merge7_split107_rready)
    ,.rresp(merge7_split107_rresp[1:0])
    ,.rvalid(merge7_split107_rvalid)
    ,.wdata(merge7_split107_wdata[(DWID - 1):0])
    ,.wlast(merge7_split107_wlast)
    ,.wready(merge7_split107_wready)
    ,.wstrb(merge7_split107_wstrb[(WSTRB - 1):0])
    ,.wvalid(merge7_split107_wvalid)

    ,.a_araddr(split107_merge210_araddr[31:0])
    ,.a_arburst(split107_merge210_arburst[1:0])
    ,.a_arextras(split107_merge210_arextras[(EXTRAS - 1):0])
    ,.a_arid(split107_merge210_arid[(IDWID - 1):0])
    ,.a_arlen(split107_merge210_arlen[7:0])
    ,.a_arready(split107_merge210_arready)
    ,.a_arvalid(split107_merge210_arvalid)
    ,.a_awaddr(split107_merge210_awaddr[31:0])
    ,.a_awburst(split107_merge210_awburst[1:0])
    ,.a_awextras(split107_merge210_awextras[(EXTRAS - 1):0])
    ,.a_awid(split107_merge210_awid[(IDWID - 1):0])
    ,.a_awlen(split107_merge210_awlen[7:0])
    ,.a_awready(split107_merge210_awready)
    ,.a_awvalid(split107_merge210_awvalid)
    ,.a_bid(split107_merge210_bid[(IDWID - 1):0])
    ,.a_bready(split107_merge210_bready)
    ,.a_bresp(split107_merge210_bresp[1:0])
    ,.a_bvalid(split107_merge210_bvalid)
    ,.a_rdata(split107_merge210_rdata[(DWID - 1):0])
    ,.a_rid(split107_merge210_rid[(IDWID - 1):0])
    ,.a_rlast(split107_merge210_rlast)
    ,.a_rready(split107_merge210_rready)
    ,.a_rresp(split107_merge210_rresp[1:0])
    ,.a_rvalid(split107_merge210_rvalid)
    ,.a_wdata(split107_merge210_wdata[(DWID - 1):0])
    ,.a_wlast(split107_merge210_wlast)
    ,.a_wready(split107_merge210_wready)
    ,.a_wstrb(split107_merge210_wstrb[(WSTRB - 1):0])
    ,.a_wvalid(split107_merge210_wvalid)
    ,.b_araddr(split107_merge202_araddr[31:0])
    ,.b_arburst(split107_merge202_arburst[1:0])
    ,.b_arextras(split107_merge202_arextras[(EXTRAS - 1):0])
    ,.b_arid(split107_merge202_arid[(IDWID - 1):0])
    ,.b_arlen(split107_merge202_arlen[7:0])
    ,.b_arready(split107_merge202_arready)
    ,.b_arvalid(split107_merge202_arvalid)
    ,.b_awaddr(split107_merge202_awaddr[31:0])
    ,.b_awburst(split107_merge202_awburst[1:0])
    ,.b_awextras(split107_merge202_awextras[(EXTRAS - 1):0])
    ,.b_awid(split107_merge202_awid[(IDWID - 1):0])
    ,.b_awlen(split107_merge202_awlen[7:0])
    ,.b_awready(split107_merge202_awready)
    ,.b_awvalid(split107_merge202_awvalid)
    ,.b_bid(split107_merge202_bid[(IDWID - 1):0])
    ,.b_bready(split107_merge202_bready)
    ,.b_bresp(split107_merge202_bresp[1:0])
    ,.b_bvalid(split107_merge202_bvalid)
    ,.b_rdata(split107_merge202_rdata[(DWID - 1):0])
    ,.b_rid(split107_merge202_rid[(IDWID - 1):0])
    ,.b_rlast(split107_merge202_rlast)
    ,.b_rready(split107_merge202_rready)
    ,.b_rresp(split107_merge202_rresp[1:0])
    ,.b_rvalid(split107_merge202_rvalid)
    ,.b_wdata(split107_merge202_wdata[(DWID - 1):0])
    ,.b_wlast(split107_merge202_wlast)
    ,.b_wready(split107_merge202_wready)
    ,.b_wstrb(split107_merge202_wstrb[(WSTRB - 1):0])
    ,.b_wvalid(split107_merge202_wvalid)
    ,.c_araddr(split107_merge207_araddr[31:0])
    ,.c_arburst(split107_merge207_arburst[1:0])
    ,.c_arextras(split107_merge207_arextras[(EXTRAS - 1):0])
    ,.c_arid(split107_merge207_arid[(IDWID - 1):0])
    ,.c_arlen(split107_merge207_arlen[7:0])
    ,.c_arready(split107_merge207_arready)
    ,.c_arvalid(split107_merge207_arvalid)
    ,.c_awaddr(split107_merge207_awaddr[31:0])
    ,.c_awburst(split107_merge207_awburst[1:0])
    ,.c_awextras(split107_merge207_awextras[(EXTRAS - 1):0])
    ,.c_awid(split107_merge207_awid[(IDWID - 1):0])
    ,.c_awlen(split107_merge207_awlen[7:0])
    ,.c_awready(split107_merge207_awready)
    ,.c_awvalid(split107_merge207_awvalid)
    ,.c_bid(split107_merge207_bid[(IDWID - 1):0])
    ,.c_bready(split107_merge207_bready)
    ,.c_bresp(split107_merge207_bresp[1:0])
    ,.c_bvalid(split107_merge207_bvalid)
    ,.c_rdata(split107_merge207_rdata[(DWID - 1):0])
    ,.c_rid(split107_merge207_rid[(IDWID - 1):0])
    ,.c_rlast(split107_merge207_rlast)
    ,.c_rready(split107_merge207_rready)
    ,.c_rresp(split107_merge207_rresp[1:0])
    ,.c_rvalid(split107_merge207_rvalid)
    ,.c_wdata(split107_merge207_wdata[(DWID - 1):0])
    ,.c_wlast(split107_merge207_wlast)
    ,.c_wready(split107_merge207_wready)
    ,.c_wstrb(split107_merge207_wstrb[(WSTRB - 1):0])
    ,.c_wvalid(split107_merge207_wvalid)
    ,.d_araddr(split107_merge211_araddr[31:0])
    ,.d_arburst(split107_merge211_arburst[1:0])
    ,.d_arextras(split107_merge211_arextras[(EXTRAS - 1):0])
    ,.d_arid(split107_merge211_arid[(IDWID - 1):0])
    ,.d_arlen(split107_merge211_arlen[7:0])
    ,.d_arready(split107_merge211_arready)
    ,.d_arvalid(split107_merge211_arvalid)
    ,.d_awaddr(split107_merge211_awaddr[31:0])
    ,.d_awburst(split107_merge211_awburst[1:0])
    ,.d_awextras(split107_merge211_awextras[(EXTRAS - 1):0])
    ,.d_awid(split107_merge211_awid[(IDWID - 1):0])
    ,.d_awlen(split107_merge211_awlen[7:0])
    ,.d_awready(split107_merge211_awready)
    ,.d_awvalid(split107_merge211_awvalid)
    ,.d_bid(split107_merge211_bid[(IDWID - 1):0])
    ,.d_bready(split107_merge211_bready)
    ,.d_bresp(split107_merge211_bresp[1:0])
    ,.d_bvalid(split107_merge211_bvalid)
    ,.d_rdata(split107_merge211_rdata[(DWID - 1):0])
    ,.d_rid(split107_merge211_rid[(IDWID - 1):0])
    ,.d_rlast(split107_merge211_rlast)
    ,.d_rready(split107_merge211_rready)
    ,.d_rresp(split107_merge211_rresp[1:0])
    ,.d_rvalid(split107_merge211_rvalid)
    ,.d_wdata(split107_merge211_wdata[(DWID - 1):0])
    ,.d_wlast(split107_merge211_wlast)
    ,.d_wready(split107_merge211_wready)
    ,.d_wstrb(split107_merge211_wstrb[(WSTRB - 1):0])
    ,.d_wvalid(split107_merge211_wvalid)

);

wire [IDWID-1:0] split108_merge211_arid ;
wire [31:0] split108_merge211_araddr ;
wire [7:0] split108_merge211_arlen ;
wire [EXTRAS-1:0] split108_merge211_arextras ;
wire [1:0] split108_merge211_arburst ;
wire split108_merge211_arvalid ;
wire split108_merge211_arready ;
wire [IDWID-1:0] split108_merge211_rid ;
wire [DWID-1:0] split108_merge211_rdata ;
wire [1:0] split108_merge211_rresp ;
wire split108_merge211_rlast ;
wire split108_merge211_rvalid ;
wire split108_merge211_rready ;

wire [IDWID-1:0] split108_merge211_awid ;
wire [31:0] split108_merge211_awaddr ;
wire [7:0] split108_merge211_awlen ;
wire [EXTRAS-1:0] split108_merge211_awextras ;
wire [1:0] split108_merge211_awburst ;
wire split108_merge211_awvalid ;
wire split108_merge211_awready ;
wire [DWID-1:0] split108_merge211_wdata ;
wire [WSTRB-1:0] split108_merge211_wstrb ;
wire split108_merge211_wlast ;
wire split108_merge211_wvalid ;
wire split108_merge211_wready ;
wire [IDWID-1:0] split108_merge211_bid ;
wire [1:0] split108_merge211_bresp ;
wire split108_merge211_bvalid ;
wire split108_merge211_bready ;


wire [IDWID-1:0] split108_merge202_arid ;
wire [31:0] split108_merge202_araddr ;
wire [7:0] split108_merge202_arlen ;
wire [EXTRAS-1:0] split108_merge202_arextras ;
wire [1:0] split108_merge202_arburst ;
wire split108_merge202_arvalid ;
wire split108_merge202_arready ;
wire [IDWID-1:0] split108_merge202_rid ;
wire [DWID-1:0] split108_merge202_rdata ;
wire [1:0] split108_merge202_rresp ;
wire split108_merge202_rlast ;
wire split108_merge202_rvalid ;
wire split108_merge202_rready ;

wire [IDWID-1:0] split108_merge202_awid ;
wire [31:0] split108_merge202_awaddr ;
wire [7:0] split108_merge202_awlen ;
wire [EXTRAS-1:0] split108_merge202_awextras ;
wire [1:0] split108_merge202_awburst ;
wire split108_merge202_awvalid ;
wire split108_merge202_awready ;
wire [DWID-1:0] split108_merge202_wdata ;
wire [WSTRB-1:0] split108_merge202_wstrb ;
wire split108_merge202_wlast ;
wire split108_merge202_wvalid ;
wire split108_merge202_wready ;
wire [IDWID-1:0] split108_merge202_bid ;
wire [1:0] split108_merge202_bresp ;
wire split108_merge202_bvalid ;
wire split108_merge202_bready ;


wire [IDWID-1:0] split108_merge205_arid ;
wire [31:0] split108_merge205_araddr ;
wire [7:0] split108_merge205_arlen ;
wire [EXTRAS-1:0] split108_merge205_arextras ;
wire [1:0] split108_merge205_arburst ;
wire split108_merge205_arvalid ;
wire split108_merge205_arready ;
wire [IDWID-1:0] split108_merge205_rid ;
wire [DWID-1:0] split108_merge205_rdata ;
wire [1:0] split108_merge205_rresp ;
wire split108_merge205_rlast ;
wire split108_merge205_rvalid ;
wire split108_merge205_rready ;

wire [IDWID-1:0] split108_merge205_awid ;
wire [31:0] split108_merge205_awaddr ;
wire [7:0] split108_merge205_awlen ;
wire [EXTRAS-1:0] split108_merge205_awextras ;
wire [1:0] split108_merge205_awburst ;
wire split108_merge205_awvalid ;
wire split108_merge205_awready ;
wire [DWID-1:0] split108_merge205_wdata ;
wire [WSTRB-1:0] split108_merge205_wstrb ;
wire split108_merge205_wlast ;
wire split108_merge205_wvalid ;
wire split108_merge205_wready ;
wire [IDWID-1:0] split108_merge205_bid ;
wire [1:0] split108_merge205_bresp ;
wire split108_merge205_bvalid ;
wire split108_merge205_bready ;


wire [IDWID-1:0] split108_merge200_arid ;
wire [31:0] split108_merge200_araddr ;
wire [7:0] split108_merge200_arlen ;
wire [EXTRAS-1:0] split108_merge200_arextras ;
wire [1:0] split108_merge200_arburst ;
wire split108_merge200_arvalid ;
wire split108_merge200_arready ;
wire [IDWID-1:0] split108_merge200_rid ;
wire [DWID-1:0] split108_merge200_rdata ;
wire [1:0] split108_merge200_rresp ;
wire split108_merge200_rlast ;
wire split108_merge200_rvalid ;
wire split108_merge200_rready ;

wire [IDWID-1:0] split108_merge200_awid ;
wire [31:0] split108_merge200_awaddr ;
wire [7:0] split108_merge200_awlen ;
wire [EXTRAS-1:0] split108_merge200_awextras ;
wire [1:0] split108_merge200_awburst ;
wire split108_merge200_awvalid ;
wire split108_merge200_awready ;
wire [DWID-1:0] split108_merge200_wdata ;
wire [WSTRB-1:0] split108_merge200_wstrb ;
wire split108_merge200_wlast ;
wire split108_merge200_wvalid ;
wire split108_merge200_wready ;
wire [IDWID-1:0] split108_merge200_bid ;
wire [1:0] split108_merge200_bresp ;
wire split108_merge200_bvalid ;
wire split108_merge200_bready ;


axi_4_splitter split108 (
     .clk(clk) ,.rst_n(rst_n)

    ,.araddr(merge8_split108_araddr[31:0])
    ,.arburst(merge8_split108_arburst[1:0])
    ,.arextras(merge8_split108_arextras[(EXTRAS - 1):0])
    ,.arid(merge8_split108_arid[(IDWID - 1):0])
    ,.arlen(merge8_split108_arlen[7:0])
    ,.arready(merge8_split108_arready)
    ,.arvalid(merge8_split108_arvalid)
    ,.awaddr(merge8_split108_awaddr[31:0])
    ,.awburst(merge8_split108_awburst[1:0])
    ,.awextras(merge8_split108_awextras[(EXTRAS - 1):0])
    ,.awid(merge8_split108_awid[3:0])
    ,.awlen(merge8_split108_awlen[7:0])
    ,.awready(merge8_split108_awready)
    ,.awvalid(merge8_split108_awvalid)
    ,.bid(merge8_split108_bid[(IDWID - 1):0])
    ,.bready(merge8_split108_bready)
    ,.bresp(merge8_split108_bresp[1:0])
    ,.bvalid(merge8_split108_bvalid)
    ,.rdata(merge8_split108_rdata[(DWID - 1):0])
    ,.rid(merge8_split108_rid[(IDWID - 1):0])
    ,.rlast(merge8_split108_rlast)
    ,.rready(merge8_split108_rready)
    ,.rresp(merge8_split108_rresp[1:0])
    ,.rvalid(merge8_split108_rvalid)
    ,.wdata(merge8_split108_wdata[(DWID - 1):0])
    ,.wlast(merge8_split108_wlast)
    ,.wready(merge8_split108_wready)
    ,.wstrb(merge8_split108_wstrb[(WSTRB - 1):0])
    ,.wvalid(merge8_split108_wvalid)

    ,.a_araddr(split108_merge211_araddr[31:0])
    ,.a_arburst(split108_merge211_arburst[1:0])
    ,.a_arextras(split108_merge211_arextras[(EXTRAS - 1):0])
    ,.a_arid(split108_merge211_arid[(IDWID - 1):0])
    ,.a_arlen(split108_merge211_arlen[7:0])
    ,.a_arready(split108_merge211_arready)
    ,.a_arvalid(split108_merge211_arvalid)
    ,.a_awaddr(split108_merge211_awaddr[31:0])
    ,.a_awburst(split108_merge211_awburst[1:0])
    ,.a_awextras(split108_merge211_awextras[(EXTRAS - 1):0])
    ,.a_awid(split108_merge211_awid[(IDWID - 1):0])
    ,.a_awlen(split108_merge211_awlen[7:0])
    ,.a_awready(split108_merge211_awready)
    ,.a_awvalid(split108_merge211_awvalid)
    ,.a_bid(split108_merge211_bid[(IDWID - 1):0])
    ,.a_bready(split108_merge211_bready)
    ,.a_bresp(split108_merge211_bresp[1:0])
    ,.a_bvalid(split108_merge211_bvalid)
    ,.a_rdata(split108_merge211_rdata[(DWID - 1):0])
    ,.a_rid(split108_merge211_rid[(IDWID - 1):0])
    ,.a_rlast(split108_merge211_rlast)
    ,.a_rready(split108_merge211_rready)
    ,.a_rresp(split108_merge211_rresp[1:0])
    ,.a_rvalid(split108_merge211_rvalid)
    ,.a_wdata(split108_merge211_wdata[(DWID - 1):0])
    ,.a_wlast(split108_merge211_wlast)
    ,.a_wready(split108_merge211_wready)
    ,.a_wstrb(split108_merge211_wstrb[(WSTRB - 1):0])
    ,.a_wvalid(split108_merge211_wvalid)
    ,.b_araddr(split108_merge202_araddr[31:0])
    ,.b_arburst(split108_merge202_arburst[1:0])
    ,.b_arextras(split108_merge202_arextras[(EXTRAS - 1):0])
    ,.b_arid(split108_merge202_arid[(IDWID - 1):0])
    ,.b_arlen(split108_merge202_arlen[7:0])
    ,.b_arready(split108_merge202_arready)
    ,.b_arvalid(split108_merge202_arvalid)
    ,.b_awaddr(split108_merge202_awaddr[31:0])
    ,.b_awburst(split108_merge202_awburst[1:0])
    ,.b_awextras(split108_merge202_awextras[(EXTRAS - 1):0])
    ,.b_awid(split108_merge202_awid[(IDWID - 1):0])
    ,.b_awlen(split108_merge202_awlen[7:0])
    ,.b_awready(split108_merge202_awready)
    ,.b_awvalid(split108_merge202_awvalid)
    ,.b_bid(split108_merge202_bid[(IDWID - 1):0])
    ,.b_bready(split108_merge202_bready)
    ,.b_bresp(split108_merge202_bresp[1:0])
    ,.b_bvalid(split108_merge202_bvalid)
    ,.b_rdata(split108_merge202_rdata[(DWID - 1):0])
    ,.b_rid(split108_merge202_rid[(IDWID - 1):0])
    ,.b_rlast(split108_merge202_rlast)
    ,.b_rready(split108_merge202_rready)
    ,.b_rresp(split108_merge202_rresp[1:0])
    ,.b_rvalid(split108_merge202_rvalid)
    ,.b_wdata(split108_merge202_wdata[(DWID - 1):0])
    ,.b_wlast(split108_merge202_wlast)
    ,.b_wready(split108_merge202_wready)
    ,.b_wstrb(split108_merge202_wstrb[(WSTRB - 1):0])
    ,.b_wvalid(split108_merge202_wvalid)
    ,.c_araddr(split108_merge205_araddr[31:0])
    ,.c_arburst(split108_merge205_arburst[1:0])
    ,.c_arextras(split108_merge205_arextras[(EXTRAS - 1):0])
    ,.c_arid(split108_merge205_arid[(IDWID - 1):0])
    ,.c_arlen(split108_merge205_arlen[7:0])
    ,.c_arready(split108_merge205_arready)
    ,.c_arvalid(split108_merge205_arvalid)
    ,.c_awaddr(split108_merge205_awaddr[31:0])
    ,.c_awburst(split108_merge205_awburst[1:0])
    ,.c_awextras(split108_merge205_awextras[(EXTRAS - 1):0])
    ,.c_awid(split108_merge205_awid[(IDWID - 1):0])
    ,.c_awlen(split108_merge205_awlen[7:0])
    ,.c_awready(split108_merge205_awready)
    ,.c_awvalid(split108_merge205_awvalid)
    ,.c_bid(split108_merge205_bid[(IDWID - 1):0])
    ,.c_bready(split108_merge205_bready)
    ,.c_bresp(split108_merge205_bresp[1:0])
    ,.c_bvalid(split108_merge205_bvalid)
    ,.c_rdata(split108_merge205_rdata[(DWID - 1):0])
    ,.c_rid(split108_merge205_rid[(IDWID - 1):0])
    ,.c_rlast(split108_merge205_rlast)
    ,.c_rready(split108_merge205_rready)
    ,.c_rresp(split108_merge205_rresp[1:0])
    ,.c_rvalid(split108_merge205_rvalid)
    ,.c_wdata(split108_merge205_wdata[(DWID - 1):0])
    ,.c_wlast(split108_merge205_wlast)
    ,.c_wready(split108_merge205_wready)
    ,.c_wstrb(split108_merge205_wstrb[(WSTRB - 1):0])
    ,.c_wvalid(split108_merge205_wvalid)
    ,.d_araddr(split108_merge200_araddr[31:0])
    ,.d_arburst(split108_merge200_arburst[1:0])
    ,.d_arextras(split108_merge200_arextras[(EXTRAS - 1):0])
    ,.d_arid(split108_merge200_arid[(IDWID - 1):0])
    ,.d_arlen(split108_merge200_arlen[7:0])
    ,.d_arready(split108_merge200_arready)
    ,.d_arvalid(split108_merge200_arvalid)
    ,.d_awaddr(split108_merge200_awaddr[31:0])
    ,.d_awburst(split108_merge200_awburst[1:0])
    ,.d_awextras(split108_merge200_awextras[(EXTRAS - 1):0])
    ,.d_awid(split108_merge200_awid[(IDWID - 1):0])
    ,.d_awlen(split108_merge200_awlen[7:0])
    ,.d_awready(split108_merge200_awready)
    ,.d_awvalid(split108_merge200_awvalid)
    ,.d_bid(split108_merge200_bid[(IDWID - 1):0])
    ,.d_bready(split108_merge200_bready)
    ,.d_bresp(split108_merge200_bresp[1:0])
    ,.d_bvalid(split108_merge200_bvalid)
    ,.d_rdata(split108_merge200_rdata[(DWID - 1):0])
    ,.d_rid(split108_merge200_rid[(IDWID - 1):0])
    ,.d_rlast(split108_merge200_rlast)
    ,.d_rready(split108_merge200_rready)
    ,.d_rresp(split108_merge200_rresp[1:0])
    ,.d_rvalid(split108_merge200_rvalid)
    ,.d_wdata(split108_merge200_wdata[(DWID - 1):0])
    ,.d_wlast(split108_merge200_wlast)
    ,.d_wready(split108_merge200_wready)
    ,.d_wstrb(split108_merge200_wstrb[(WSTRB - 1):0])
    ,.d_wvalid(split108_merge200_wvalid)

);

wire [IDWID-1:0] split109_merge215_arid ;
wire [31:0] split109_merge215_araddr ;
wire [7:0] split109_merge215_arlen ;
wire [EXTRAS-1:0] split109_merge215_arextras ;
wire [1:0] split109_merge215_arburst ;
wire split109_merge215_arvalid ;
wire split109_merge215_arready ;
wire [IDWID-1:0] split109_merge215_rid ;
wire [DWID-1:0] split109_merge215_rdata ;
wire [1:0] split109_merge215_rresp ;
wire split109_merge215_rlast ;
wire split109_merge215_rvalid ;
wire split109_merge215_rready ;

wire [IDWID-1:0] split109_merge215_awid ;
wire [31:0] split109_merge215_awaddr ;
wire [7:0] split109_merge215_awlen ;
wire [EXTRAS-1:0] split109_merge215_awextras ;
wire [1:0] split109_merge215_awburst ;
wire split109_merge215_awvalid ;
wire split109_merge215_awready ;
wire [DWID-1:0] split109_merge215_wdata ;
wire [WSTRB-1:0] split109_merge215_wstrb ;
wire split109_merge215_wlast ;
wire split109_merge215_wvalid ;
wire split109_merge215_wready ;
wire [IDWID-1:0] split109_merge215_bid ;
wire [1:0] split109_merge215_bresp ;
wire split109_merge215_bvalid ;
wire split109_merge215_bready ;


wire [IDWID-1:0] split109_merge209_arid ;
wire [31:0] split109_merge209_araddr ;
wire [7:0] split109_merge209_arlen ;
wire [EXTRAS-1:0] split109_merge209_arextras ;
wire [1:0] split109_merge209_arburst ;
wire split109_merge209_arvalid ;
wire split109_merge209_arready ;
wire [IDWID-1:0] split109_merge209_rid ;
wire [DWID-1:0] split109_merge209_rdata ;
wire [1:0] split109_merge209_rresp ;
wire split109_merge209_rlast ;
wire split109_merge209_rvalid ;
wire split109_merge209_rready ;

wire [IDWID-1:0] split109_merge209_awid ;
wire [31:0] split109_merge209_awaddr ;
wire [7:0] split109_merge209_awlen ;
wire [EXTRAS-1:0] split109_merge209_awextras ;
wire [1:0] split109_merge209_awburst ;
wire split109_merge209_awvalid ;
wire split109_merge209_awready ;
wire [DWID-1:0] split109_merge209_wdata ;
wire [WSTRB-1:0] split109_merge209_wstrb ;
wire split109_merge209_wlast ;
wire split109_merge209_wvalid ;
wire split109_merge209_wready ;
wire [IDWID-1:0] split109_merge209_bid ;
wire [1:0] split109_merge209_bresp ;
wire split109_merge209_bvalid ;
wire split109_merge209_bready ;


wire [IDWID-1:0] split109_merge204_arid ;
wire [31:0] split109_merge204_araddr ;
wire [7:0] split109_merge204_arlen ;
wire [EXTRAS-1:0] split109_merge204_arextras ;
wire [1:0] split109_merge204_arburst ;
wire split109_merge204_arvalid ;
wire split109_merge204_arready ;
wire [IDWID-1:0] split109_merge204_rid ;
wire [DWID-1:0] split109_merge204_rdata ;
wire [1:0] split109_merge204_rresp ;
wire split109_merge204_rlast ;
wire split109_merge204_rvalid ;
wire split109_merge204_rready ;

wire [IDWID-1:0] split109_merge204_awid ;
wire [31:0] split109_merge204_awaddr ;
wire [7:0] split109_merge204_awlen ;
wire [EXTRAS-1:0] split109_merge204_awextras ;
wire [1:0] split109_merge204_awburst ;
wire split109_merge204_awvalid ;
wire split109_merge204_awready ;
wire [DWID-1:0] split109_merge204_wdata ;
wire [WSTRB-1:0] split109_merge204_wstrb ;
wire split109_merge204_wlast ;
wire split109_merge204_wvalid ;
wire split109_merge204_wready ;
wire [IDWID-1:0] split109_merge204_bid ;
wire [1:0] split109_merge204_bresp ;
wire split109_merge204_bvalid ;
wire split109_merge204_bready ;


wire [IDWID-1:0] split109_merge203_arid ;
wire [31:0] split109_merge203_araddr ;
wire [7:0] split109_merge203_arlen ;
wire [EXTRAS-1:0] split109_merge203_arextras ;
wire [1:0] split109_merge203_arburst ;
wire split109_merge203_arvalid ;
wire split109_merge203_arready ;
wire [IDWID-1:0] split109_merge203_rid ;
wire [DWID-1:0] split109_merge203_rdata ;
wire [1:0] split109_merge203_rresp ;
wire split109_merge203_rlast ;
wire split109_merge203_rvalid ;
wire split109_merge203_rready ;

wire [IDWID-1:0] split109_merge203_awid ;
wire [31:0] split109_merge203_awaddr ;
wire [7:0] split109_merge203_awlen ;
wire [EXTRAS-1:0] split109_merge203_awextras ;
wire [1:0] split109_merge203_awburst ;
wire split109_merge203_awvalid ;
wire split109_merge203_awready ;
wire [DWID-1:0] split109_merge203_wdata ;
wire [WSTRB-1:0] split109_merge203_wstrb ;
wire split109_merge203_wlast ;
wire split109_merge203_wvalid ;
wire split109_merge203_wready ;
wire [IDWID-1:0] split109_merge203_bid ;
wire [1:0] split109_merge203_bresp ;
wire split109_merge203_bvalid ;
wire split109_merge203_bready ;


axi_4_splitter split109 (
     .clk(clk) ,.rst_n(rst_n)

    ,.araddr(merge9_split109_araddr[31:0])
    ,.arburst(merge9_split109_arburst[1:0])
    ,.arextras(merge9_split109_arextras[(EXTRAS - 1):0])
    ,.arid(merge9_split109_arid[(IDWID - 1):0])
    ,.arlen(merge9_split109_arlen[7:0])
    ,.arready(merge9_split109_arready)
    ,.arvalid(merge9_split109_arvalid)
    ,.awaddr(merge9_split109_awaddr[31:0])
    ,.awburst(merge9_split109_awburst[1:0])
    ,.awextras(merge9_split109_awextras[(EXTRAS - 1):0])
    ,.awid(merge9_split109_awid[3:0])
    ,.awlen(merge9_split109_awlen[7:0])
    ,.awready(merge9_split109_awready)
    ,.awvalid(merge9_split109_awvalid)
    ,.bid(merge9_split109_bid[(IDWID - 1):0])
    ,.bready(merge9_split109_bready)
    ,.bresp(merge9_split109_bresp[1:0])
    ,.bvalid(merge9_split109_bvalid)
    ,.rdata(merge9_split109_rdata[(DWID - 1):0])
    ,.rid(merge9_split109_rid[(IDWID - 1):0])
    ,.rlast(merge9_split109_rlast)
    ,.rready(merge9_split109_rready)
    ,.rresp(merge9_split109_rresp[1:0])
    ,.rvalid(merge9_split109_rvalid)
    ,.wdata(merge9_split109_wdata[(DWID - 1):0])
    ,.wlast(merge9_split109_wlast)
    ,.wready(merge9_split109_wready)
    ,.wstrb(merge9_split109_wstrb[(WSTRB - 1):0])
    ,.wvalid(merge9_split109_wvalid)

    ,.a_araddr(split109_merge215_araddr[31:0])
    ,.a_arburst(split109_merge215_arburst[1:0])
    ,.a_arextras(split109_merge215_arextras[(EXTRAS - 1):0])
    ,.a_arid(split109_merge215_arid[(IDWID - 1):0])
    ,.a_arlen(split109_merge215_arlen[7:0])
    ,.a_arready(split109_merge215_arready)
    ,.a_arvalid(split109_merge215_arvalid)
    ,.a_awaddr(split109_merge215_awaddr[31:0])
    ,.a_awburst(split109_merge215_awburst[1:0])
    ,.a_awextras(split109_merge215_awextras[(EXTRAS - 1):0])
    ,.a_awid(split109_merge215_awid[(IDWID - 1):0])
    ,.a_awlen(split109_merge215_awlen[7:0])
    ,.a_awready(split109_merge215_awready)
    ,.a_awvalid(split109_merge215_awvalid)
    ,.a_bid(split109_merge215_bid[(IDWID - 1):0])
    ,.a_bready(split109_merge215_bready)
    ,.a_bresp(split109_merge215_bresp[1:0])
    ,.a_bvalid(split109_merge215_bvalid)
    ,.a_rdata(split109_merge215_rdata[(DWID - 1):0])
    ,.a_rid(split109_merge215_rid[(IDWID - 1):0])
    ,.a_rlast(split109_merge215_rlast)
    ,.a_rready(split109_merge215_rready)
    ,.a_rresp(split109_merge215_rresp[1:0])
    ,.a_rvalid(split109_merge215_rvalid)
    ,.a_wdata(split109_merge215_wdata[(DWID - 1):0])
    ,.a_wlast(split109_merge215_wlast)
    ,.a_wready(split109_merge215_wready)
    ,.a_wstrb(split109_merge215_wstrb[(WSTRB - 1):0])
    ,.a_wvalid(split109_merge215_wvalid)
    ,.b_araddr(split109_merge209_araddr[31:0])
    ,.b_arburst(split109_merge209_arburst[1:0])
    ,.b_arextras(split109_merge209_arextras[(EXTRAS - 1):0])
    ,.b_arid(split109_merge209_arid[(IDWID - 1):0])
    ,.b_arlen(split109_merge209_arlen[7:0])
    ,.b_arready(split109_merge209_arready)
    ,.b_arvalid(split109_merge209_arvalid)
    ,.b_awaddr(split109_merge209_awaddr[31:0])
    ,.b_awburst(split109_merge209_awburst[1:0])
    ,.b_awextras(split109_merge209_awextras[(EXTRAS - 1):0])
    ,.b_awid(split109_merge209_awid[(IDWID - 1):0])
    ,.b_awlen(split109_merge209_awlen[7:0])
    ,.b_awready(split109_merge209_awready)
    ,.b_awvalid(split109_merge209_awvalid)
    ,.b_bid(split109_merge209_bid[(IDWID - 1):0])
    ,.b_bready(split109_merge209_bready)
    ,.b_bresp(split109_merge209_bresp[1:0])
    ,.b_bvalid(split109_merge209_bvalid)
    ,.b_rdata(split109_merge209_rdata[(DWID - 1):0])
    ,.b_rid(split109_merge209_rid[(IDWID - 1):0])
    ,.b_rlast(split109_merge209_rlast)
    ,.b_rready(split109_merge209_rready)
    ,.b_rresp(split109_merge209_rresp[1:0])
    ,.b_rvalid(split109_merge209_rvalid)
    ,.b_wdata(split109_merge209_wdata[(DWID - 1):0])
    ,.b_wlast(split109_merge209_wlast)
    ,.b_wready(split109_merge209_wready)
    ,.b_wstrb(split109_merge209_wstrb[(WSTRB - 1):0])
    ,.b_wvalid(split109_merge209_wvalid)
    ,.c_araddr(split109_merge204_araddr[31:0])
    ,.c_arburst(split109_merge204_arburst[1:0])
    ,.c_arextras(split109_merge204_arextras[(EXTRAS - 1):0])
    ,.c_arid(split109_merge204_arid[(IDWID - 1):0])
    ,.c_arlen(split109_merge204_arlen[7:0])
    ,.c_arready(split109_merge204_arready)
    ,.c_arvalid(split109_merge204_arvalid)
    ,.c_awaddr(split109_merge204_awaddr[31:0])
    ,.c_awburst(split109_merge204_awburst[1:0])
    ,.c_awextras(split109_merge204_awextras[(EXTRAS - 1):0])
    ,.c_awid(split109_merge204_awid[(IDWID - 1):0])
    ,.c_awlen(split109_merge204_awlen[7:0])
    ,.c_awready(split109_merge204_awready)
    ,.c_awvalid(split109_merge204_awvalid)
    ,.c_bid(split109_merge204_bid[(IDWID - 1):0])
    ,.c_bready(split109_merge204_bready)
    ,.c_bresp(split109_merge204_bresp[1:0])
    ,.c_bvalid(split109_merge204_bvalid)
    ,.c_rdata(split109_merge204_rdata[(DWID - 1):0])
    ,.c_rid(split109_merge204_rid[(IDWID - 1):0])
    ,.c_rlast(split109_merge204_rlast)
    ,.c_rready(split109_merge204_rready)
    ,.c_rresp(split109_merge204_rresp[1:0])
    ,.c_rvalid(split109_merge204_rvalid)
    ,.c_wdata(split109_merge204_wdata[(DWID - 1):0])
    ,.c_wlast(split109_merge204_wlast)
    ,.c_wready(split109_merge204_wready)
    ,.c_wstrb(split109_merge204_wstrb[(WSTRB - 1):0])
    ,.c_wvalid(split109_merge204_wvalid)
    ,.d_araddr(split109_merge203_araddr[31:0])
    ,.d_arburst(split109_merge203_arburst[1:0])
    ,.d_arextras(split109_merge203_arextras[(EXTRAS - 1):0])
    ,.d_arid(split109_merge203_arid[(IDWID - 1):0])
    ,.d_arlen(split109_merge203_arlen[7:0])
    ,.d_arready(split109_merge203_arready)
    ,.d_arvalid(split109_merge203_arvalid)
    ,.d_awaddr(split109_merge203_awaddr[31:0])
    ,.d_awburst(split109_merge203_awburst[1:0])
    ,.d_awextras(split109_merge203_awextras[(EXTRAS - 1):0])
    ,.d_awid(split109_merge203_awid[(IDWID - 1):0])
    ,.d_awlen(split109_merge203_awlen[7:0])
    ,.d_awready(split109_merge203_awready)
    ,.d_awvalid(split109_merge203_awvalid)
    ,.d_bid(split109_merge203_bid[(IDWID - 1):0])
    ,.d_bready(split109_merge203_bready)
    ,.d_bresp(split109_merge203_bresp[1:0])
    ,.d_bvalid(split109_merge203_bvalid)
    ,.d_rdata(split109_merge203_rdata[(DWID - 1):0])
    ,.d_rid(split109_merge203_rid[(IDWID - 1):0])
    ,.d_rlast(split109_merge203_rlast)
    ,.d_rready(split109_merge203_rready)
    ,.d_rresp(split109_merge203_rresp[1:0])
    ,.d_rvalid(split109_merge203_rvalid)
    ,.d_wdata(split109_merge203_wdata[(DWID - 1):0])
    ,.d_wlast(split109_merge203_wlast)
    ,.d_wready(split109_merge203_wready)
    ,.d_wstrb(split109_merge203_wstrb[(WSTRB - 1):0])
    ,.d_wvalid(split109_merge203_wvalid)

);

wire [IDWID-1:0] split110_merge215_arid ;
wire [31:0] split110_merge215_araddr ;
wire [7:0] split110_merge215_arlen ;
wire [EXTRAS-1:0] split110_merge215_arextras ;
wire [1:0] split110_merge215_arburst ;
wire split110_merge215_arvalid ;
wire split110_merge215_arready ;
wire [IDWID-1:0] split110_merge215_rid ;
wire [DWID-1:0] split110_merge215_rdata ;
wire [1:0] split110_merge215_rresp ;
wire split110_merge215_rlast ;
wire split110_merge215_rvalid ;
wire split110_merge215_rready ;

wire [IDWID-1:0] split110_merge215_awid ;
wire [31:0] split110_merge215_awaddr ;
wire [7:0] split110_merge215_awlen ;
wire [EXTRAS-1:0] split110_merge215_awextras ;
wire [1:0] split110_merge215_awburst ;
wire split110_merge215_awvalid ;
wire split110_merge215_awready ;
wire [DWID-1:0] split110_merge215_wdata ;
wire [WSTRB-1:0] split110_merge215_wstrb ;
wire split110_merge215_wlast ;
wire split110_merge215_wvalid ;
wire split110_merge215_wready ;
wire [IDWID-1:0] split110_merge215_bid ;
wire [1:0] split110_merge215_bresp ;
wire split110_merge215_bvalid ;
wire split110_merge215_bready ;


wire [IDWID-1:0] split110_merge203_arid ;
wire [31:0] split110_merge203_araddr ;
wire [7:0] split110_merge203_arlen ;
wire [EXTRAS-1:0] split110_merge203_arextras ;
wire [1:0] split110_merge203_arburst ;
wire split110_merge203_arvalid ;
wire split110_merge203_arready ;
wire [IDWID-1:0] split110_merge203_rid ;
wire [DWID-1:0] split110_merge203_rdata ;
wire [1:0] split110_merge203_rresp ;
wire split110_merge203_rlast ;
wire split110_merge203_rvalid ;
wire split110_merge203_rready ;

wire [IDWID-1:0] split110_merge203_awid ;
wire [31:0] split110_merge203_awaddr ;
wire [7:0] split110_merge203_awlen ;
wire [EXTRAS-1:0] split110_merge203_awextras ;
wire [1:0] split110_merge203_awburst ;
wire split110_merge203_awvalid ;
wire split110_merge203_awready ;
wire [DWID-1:0] split110_merge203_wdata ;
wire [WSTRB-1:0] split110_merge203_wstrb ;
wire split110_merge203_wlast ;
wire split110_merge203_wvalid ;
wire split110_merge203_wready ;
wire [IDWID-1:0] split110_merge203_bid ;
wire [1:0] split110_merge203_bresp ;
wire split110_merge203_bvalid ;
wire split110_merge203_bready ;


wire [IDWID-1:0] split110_merge209_arid ;
wire [31:0] split110_merge209_araddr ;
wire [7:0] split110_merge209_arlen ;
wire [EXTRAS-1:0] split110_merge209_arextras ;
wire [1:0] split110_merge209_arburst ;
wire split110_merge209_arvalid ;
wire split110_merge209_arready ;
wire [IDWID-1:0] split110_merge209_rid ;
wire [DWID-1:0] split110_merge209_rdata ;
wire [1:0] split110_merge209_rresp ;
wire split110_merge209_rlast ;
wire split110_merge209_rvalid ;
wire split110_merge209_rready ;

wire [IDWID-1:0] split110_merge209_awid ;
wire [31:0] split110_merge209_awaddr ;
wire [7:0] split110_merge209_awlen ;
wire [EXTRAS-1:0] split110_merge209_awextras ;
wire [1:0] split110_merge209_awburst ;
wire split110_merge209_awvalid ;
wire split110_merge209_awready ;
wire [DWID-1:0] split110_merge209_wdata ;
wire [WSTRB-1:0] split110_merge209_wstrb ;
wire split110_merge209_wlast ;
wire split110_merge209_wvalid ;
wire split110_merge209_wready ;
wire [IDWID-1:0] split110_merge209_bid ;
wire [1:0] split110_merge209_bresp ;
wire split110_merge209_bvalid ;
wire split110_merge209_bready ;


wire [IDWID-1:0] split110_merge214_arid ;
wire [31:0] split110_merge214_araddr ;
wire [7:0] split110_merge214_arlen ;
wire [EXTRAS-1:0] split110_merge214_arextras ;
wire [1:0] split110_merge214_arburst ;
wire split110_merge214_arvalid ;
wire split110_merge214_arready ;
wire [IDWID-1:0] split110_merge214_rid ;
wire [DWID-1:0] split110_merge214_rdata ;
wire [1:0] split110_merge214_rresp ;
wire split110_merge214_rlast ;
wire split110_merge214_rvalid ;
wire split110_merge214_rready ;

wire [IDWID-1:0] split110_merge214_awid ;
wire [31:0] split110_merge214_awaddr ;
wire [7:0] split110_merge214_awlen ;
wire [EXTRAS-1:0] split110_merge214_awextras ;
wire [1:0] split110_merge214_awburst ;
wire split110_merge214_awvalid ;
wire split110_merge214_awready ;
wire [DWID-1:0] split110_merge214_wdata ;
wire [WSTRB-1:0] split110_merge214_wstrb ;
wire split110_merge214_wlast ;
wire split110_merge214_wvalid ;
wire split110_merge214_wready ;
wire [IDWID-1:0] split110_merge214_bid ;
wire [1:0] split110_merge214_bresp ;
wire split110_merge214_bvalid ;
wire split110_merge214_bready ;


axi_4_splitter split110 (
     .clk(clk) ,.rst_n(rst_n)

    ,.araddr(merge10_split110_araddr[31:0])
    ,.arburst(merge10_split110_arburst[1:0])
    ,.arextras(merge10_split110_arextras[(EXTRAS - 1):0])
    ,.arid(merge10_split110_arid[(IDWID - 1):0])
    ,.arlen(merge10_split110_arlen[7:0])
    ,.arready(merge10_split110_arready)
    ,.arvalid(merge10_split110_arvalid)
    ,.awaddr(merge10_split110_awaddr[31:0])
    ,.awburst(merge10_split110_awburst[1:0])
    ,.awextras(merge10_split110_awextras[(EXTRAS - 1):0])
    ,.awid(merge10_split110_awid[3:0])
    ,.awlen(merge10_split110_awlen[7:0])
    ,.awready(merge10_split110_awready)
    ,.awvalid(merge10_split110_awvalid)
    ,.bid(merge10_split110_bid[(IDWID - 1):0])
    ,.bready(merge10_split110_bready)
    ,.bresp(merge10_split110_bresp[1:0])
    ,.bvalid(merge10_split110_bvalid)
    ,.rdata(merge10_split110_rdata[(DWID - 1):0])
    ,.rid(merge10_split110_rid[(IDWID - 1):0])
    ,.rlast(merge10_split110_rlast)
    ,.rready(merge10_split110_rready)
    ,.rresp(merge10_split110_rresp[1:0])
    ,.rvalid(merge10_split110_rvalid)
    ,.wdata(merge10_split110_wdata[(DWID - 1):0])
    ,.wlast(merge10_split110_wlast)
    ,.wready(merge10_split110_wready)
    ,.wstrb(merge10_split110_wstrb[(WSTRB - 1):0])
    ,.wvalid(merge10_split110_wvalid)

    ,.a_araddr(split110_merge215_araddr[31:0])
    ,.a_arburst(split110_merge215_arburst[1:0])
    ,.a_arextras(split110_merge215_arextras[(EXTRAS - 1):0])
    ,.a_arid(split110_merge215_arid[(IDWID - 1):0])
    ,.a_arlen(split110_merge215_arlen[7:0])
    ,.a_arready(split110_merge215_arready)
    ,.a_arvalid(split110_merge215_arvalid)
    ,.a_awaddr(split110_merge215_awaddr[31:0])
    ,.a_awburst(split110_merge215_awburst[1:0])
    ,.a_awextras(split110_merge215_awextras[(EXTRAS - 1):0])
    ,.a_awid(split110_merge215_awid[(IDWID - 1):0])
    ,.a_awlen(split110_merge215_awlen[7:0])
    ,.a_awready(split110_merge215_awready)
    ,.a_awvalid(split110_merge215_awvalid)
    ,.a_bid(split110_merge215_bid[(IDWID - 1):0])
    ,.a_bready(split110_merge215_bready)
    ,.a_bresp(split110_merge215_bresp[1:0])
    ,.a_bvalid(split110_merge215_bvalid)
    ,.a_rdata(split110_merge215_rdata[(DWID - 1):0])
    ,.a_rid(split110_merge215_rid[(IDWID - 1):0])
    ,.a_rlast(split110_merge215_rlast)
    ,.a_rready(split110_merge215_rready)
    ,.a_rresp(split110_merge215_rresp[1:0])
    ,.a_rvalid(split110_merge215_rvalid)
    ,.a_wdata(split110_merge215_wdata[(DWID - 1):0])
    ,.a_wlast(split110_merge215_wlast)
    ,.a_wready(split110_merge215_wready)
    ,.a_wstrb(split110_merge215_wstrb[(WSTRB - 1):0])
    ,.a_wvalid(split110_merge215_wvalid)
    ,.b_araddr(split110_merge203_araddr[31:0])
    ,.b_arburst(split110_merge203_arburst[1:0])
    ,.b_arextras(split110_merge203_arextras[(EXTRAS - 1):0])
    ,.b_arid(split110_merge203_arid[(IDWID - 1):0])
    ,.b_arlen(split110_merge203_arlen[7:0])
    ,.b_arready(split110_merge203_arready)
    ,.b_arvalid(split110_merge203_arvalid)
    ,.b_awaddr(split110_merge203_awaddr[31:0])
    ,.b_awburst(split110_merge203_awburst[1:0])
    ,.b_awextras(split110_merge203_awextras[(EXTRAS - 1):0])
    ,.b_awid(split110_merge203_awid[(IDWID - 1):0])
    ,.b_awlen(split110_merge203_awlen[7:0])
    ,.b_awready(split110_merge203_awready)
    ,.b_awvalid(split110_merge203_awvalid)
    ,.b_bid(split110_merge203_bid[(IDWID - 1):0])
    ,.b_bready(split110_merge203_bready)
    ,.b_bresp(split110_merge203_bresp[1:0])
    ,.b_bvalid(split110_merge203_bvalid)
    ,.b_rdata(split110_merge203_rdata[(DWID - 1):0])
    ,.b_rid(split110_merge203_rid[(IDWID - 1):0])
    ,.b_rlast(split110_merge203_rlast)
    ,.b_rready(split110_merge203_rready)
    ,.b_rresp(split110_merge203_rresp[1:0])
    ,.b_rvalid(split110_merge203_rvalid)
    ,.b_wdata(split110_merge203_wdata[(DWID - 1):0])
    ,.b_wlast(split110_merge203_wlast)
    ,.b_wready(split110_merge203_wready)
    ,.b_wstrb(split110_merge203_wstrb[(WSTRB - 1):0])
    ,.b_wvalid(split110_merge203_wvalid)
    ,.c_araddr(split110_merge209_araddr[31:0])
    ,.c_arburst(split110_merge209_arburst[1:0])
    ,.c_arextras(split110_merge209_arextras[(EXTRAS - 1):0])
    ,.c_arid(split110_merge209_arid[(IDWID - 1):0])
    ,.c_arlen(split110_merge209_arlen[7:0])
    ,.c_arready(split110_merge209_arready)
    ,.c_arvalid(split110_merge209_arvalid)
    ,.c_awaddr(split110_merge209_awaddr[31:0])
    ,.c_awburst(split110_merge209_awburst[1:0])
    ,.c_awextras(split110_merge209_awextras[(EXTRAS - 1):0])
    ,.c_awid(split110_merge209_awid[(IDWID - 1):0])
    ,.c_awlen(split110_merge209_awlen[7:0])
    ,.c_awready(split110_merge209_awready)
    ,.c_awvalid(split110_merge209_awvalid)
    ,.c_bid(split110_merge209_bid[(IDWID - 1):0])
    ,.c_bready(split110_merge209_bready)
    ,.c_bresp(split110_merge209_bresp[1:0])
    ,.c_bvalid(split110_merge209_bvalid)
    ,.c_rdata(split110_merge209_rdata[(DWID - 1):0])
    ,.c_rid(split110_merge209_rid[(IDWID - 1):0])
    ,.c_rlast(split110_merge209_rlast)
    ,.c_rready(split110_merge209_rready)
    ,.c_rresp(split110_merge209_rresp[1:0])
    ,.c_rvalid(split110_merge209_rvalid)
    ,.c_wdata(split110_merge209_wdata[(DWID - 1):0])
    ,.c_wlast(split110_merge209_wlast)
    ,.c_wready(split110_merge209_wready)
    ,.c_wstrb(split110_merge209_wstrb[(WSTRB - 1):0])
    ,.c_wvalid(split110_merge209_wvalid)
    ,.d_araddr(split110_merge214_araddr[31:0])
    ,.d_arburst(split110_merge214_arburst[1:0])
    ,.d_arextras(split110_merge214_arextras[(EXTRAS - 1):0])
    ,.d_arid(split110_merge214_arid[(IDWID - 1):0])
    ,.d_arlen(split110_merge214_arlen[7:0])
    ,.d_arready(split110_merge214_arready)
    ,.d_arvalid(split110_merge214_arvalid)
    ,.d_awaddr(split110_merge214_awaddr[31:0])
    ,.d_awburst(split110_merge214_awburst[1:0])
    ,.d_awextras(split110_merge214_awextras[(EXTRAS - 1):0])
    ,.d_awid(split110_merge214_awid[(IDWID - 1):0])
    ,.d_awlen(split110_merge214_awlen[7:0])
    ,.d_awready(split110_merge214_awready)
    ,.d_awvalid(split110_merge214_awvalid)
    ,.d_bid(split110_merge214_bid[(IDWID - 1):0])
    ,.d_bready(split110_merge214_bready)
    ,.d_bresp(split110_merge214_bresp[1:0])
    ,.d_bvalid(split110_merge214_bvalid)
    ,.d_rdata(split110_merge214_rdata[(DWID - 1):0])
    ,.d_rid(split110_merge214_rid[(IDWID - 1):0])
    ,.d_rlast(split110_merge214_rlast)
    ,.d_rready(split110_merge214_rready)
    ,.d_rresp(split110_merge214_rresp[1:0])
    ,.d_rvalid(split110_merge214_rvalid)
    ,.d_wdata(split110_merge214_wdata[(DWID - 1):0])
    ,.d_wlast(split110_merge214_wlast)
    ,.d_wready(split110_merge214_wready)
    ,.d_wstrb(split110_merge214_wstrb[(WSTRB - 1):0])
    ,.d_wvalid(split110_merge214_wvalid)

);

wire [IDWID-1:0] split111_merge213_arid ;
wire [31:0] split111_merge213_araddr ;
wire [7:0] split111_merge213_arlen ;
wire [EXTRAS-1:0] split111_merge213_arextras ;
wire [1:0] split111_merge213_arburst ;
wire split111_merge213_arvalid ;
wire split111_merge213_arready ;
wire [IDWID-1:0] split111_merge213_rid ;
wire [DWID-1:0] split111_merge213_rdata ;
wire [1:0] split111_merge213_rresp ;
wire split111_merge213_rlast ;
wire split111_merge213_rvalid ;
wire split111_merge213_rready ;

wire [IDWID-1:0] split111_merge213_awid ;
wire [31:0] split111_merge213_awaddr ;
wire [7:0] split111_merge213_awlen ;
wire [EXTRAS-1:0] split111_merge213_awextras ;
wire [1:0] split111_merge213_awburst ;
wire split111_merge213_awvalid ;
wire split111_merge213_awready ;
wire [DWID-1:0] split111_merge213_wdata ;
wire [WSTRB-1:0] split111_merge213_wstrb ;
wire split111_merge213_wlast ;
wire split111_merge213_wvalid ;
wire split111_merge213_wready ;
wire [IDWID-1:0] split111_merge213_bid ;
wire [1:0] split111_merge213_bresp ;
wire split111_merge213_bvalid ;
wire split111_merge213_bready ;


wire [IDWID-1:0] split111_merge200_arid ;
wire [31:0] split111_merge200_araddr ;
wire [7:0] split111_merge200_arlen ;
wire [EXTRAS-1:0] split111_merge200_arextras ;
wire [1:0] split111_merge200_arburst ;
wire split111_merge200_arvalid ;
wire split111_merge200_arready ;
wire [IDWID-1:0] split111_merge200_rid ;
wire [DWID-1:0] split111_merge200_rdata ;
wire [1:0] split111_merge200_rresp ;
wire split111_merge200_rlast ;
wire split111_merge200_rvalid ;
wire split111_merge200_rready ;

wire [IDWID-1:0] split111_merge200_awid ;
wire [31:0] split111_merge200_awaddr ;
wire [7:0] split111_merge200_awlen ;
wire [EXTRAS-1:0] split111_merge200_awextras ;
wire [1:0] split111_merge200_awburst ;
wire split111_merge200_awvalid ;
wire split111_merge200_awready ;
wire [DWID-1:0] split111_merge200_wdata ;
wire [WSTRB-1:0] split111_merge200_wstrb ;
wire split111_merge200_wlast ;
wire split111_merge200_wvalid ;
wire split111_merge200_wready ;
wire [IDWID-1:0] split111_merge200_bid ;
wire [1:0] split111_merge200_bresp ;
wire split111_merge200_bvalid ;
wire split111_merge200_bready ;


wire [IDWID-1:0] split111_merge202_arid ;
wire [31:0] split111_merge202_araddr ;
wire [7:0] split111_merge202_arlen ;
wire [EXTRAS-1:0] split111_merge202_arextras ;
wire [1:0] split111_merge202_arburst ;
wire split111_merge202_arvalid ;
wire split111_merge202_arready ;
wire [IDWID-1:0] split111_merge202_rid ;
wire [DWID-1:0] split111_merge202_rdata ;
wire [1:0] split111_merge202_rresp ;
wire split111_merge202_rlast ;
wire split111_merge202_rvalid ;
wire split111_merge202_rready ;

wire [IDWID-1:0] split111_merge202_awid ;
wire [31:0] split111_merge202_awaddr ;
wire [7:0] split111_merge202_awlen ;
wire [EXTRAS-1:0] split111_merge202_awextras ;
wire [1:0] split111_merge202_awburst ;
wire split111_merge202_awvalid ;
wire split111_merge202_awready ;
wire [DWID-1:0] split111_merge202_wdata ;
wire [WSTRB-1:0] split111_merge202_wstrb ;
wire split111_merge202_wlast ;
wire split111_merge202_wvalid ;
wire split111_merge202_wready ;
wire [IDWID-1:0] split111_merge202_bid ;
wire [1:0] split111_merge202_bresp ;
wire split111_merge202_bvalid ;
wire split111_merge202_bready ;


wire [IDWID-1:0] split111_merge214_arid ;
wire [31:0] split111_merge214_araddr ;
wire [7:0] split111_merge214_arlen ;
wire [EXTRAS-1:0] split111_merge214_arextras ;
wire [1:0] split111_merge214_arburst ;
wire split111_merge214_arvalid ;
wire split111_merge214_arready ;
wire [IDWID-1:0] split111_merge214_rid ;
wire [DWID-1:0] split111_merge214_rdata ;
wire [1:0] split111_merge214_rresp ;
wire split111_merge214_rlast ;
wire split111_merge214_rvalid ;
wire split111_merge214_rready ;

wire [IDWID-1:0] split111_merge214_awid ;
wire [31:0] split111_merge214_awaddr ;
wire [7:0] split111_merge214_awlen ;
wire [EXTRAS-1:0] split111_merge214_awextras ;
wire [1:0] split111_merge214_awburst ;
wire split111_merge214_awvalid ;
wire split111_merge214_awready ;
wire [DWID-1:0] split111_merge214_wdata ;
wire [WSTRB-1:0] split111_merge214_wstrb ;
wire split111_merge214_wlast ;
wire split111_merge214_wvalid ;
wire split111_merge214_wready ;
wire [IDWID-1:0] split111_merge214_bid ;
wire [1:0] split111_merge214_bresp ;
wire split111_merge214_bvalid ;
wire split111_merge214_bready ;


axi_4_splitter split111 (
     .clk(clk) ,.rst_n(rst_n)

    ,.araddr(merge11_split111_araddr[31:0])
    ,.arburst(merge11_split111_arburst[1:0])
    ,.arextras(merge11_split111_arextras[(EXTRAS - 1):0])
    ,.arid(merge11_split111_arid[(IDWID - 1):0])
    ,.arlen(merge11_split111_arlen[7:0])
    ,.arready(merge11_split111_arready)
    ,.arvalid(merge11_split111_arvalid)
    ,.awaddr(merge11_split111_awaddr[31:0])
    ,.awburst(merge11_split111_awburst[1:0])
    ,.awextras(merge11_split111_awextras[(EXTRAS - 1):0])
    ,.awid(merge11_split111_awid[3:0])
    ,.awlen(merge11_split111_awlen[7:0])
    ,.awready(merge11_split111_awready)
    ,.awvalid(merge11_split111_awvalid)
    ,.bid(merge11_split111_bid[(IDWID - 1):0])
    ,.bready(merge11_split111_bready)
    ,.bresp(merge11_split111_bresp[1:0])
    ,.bvalid(merge11_split111_bvalid)
    ,.rdata(merge11_split111_rdata[(DWID - 1):0])
    ,.rid(merge11_split111_rid[(IDWID - 1):0])
    ,.rlast(merge11_split111_rlast)
    ,.rready(merge11_split111_rready)
    ,.rresp(merge11_split111_rresp[1:0])
    ,.rvalid(merge11_split111_rvalid)
    ,.wdata(merge11_split111_wdata[(DWID - 1):0])
    ,.wlast(merge11_split111_wlast)
    ,.wready(merge11_split111_wready)
    ,.wstrb(merge11_split111_wstrb[(WSTRB - 1):0])
    ,.wvalid(merge11_split111_wvalid)

    ,.a_araddr(split111_merge213_araddr[31:0])
    ,.a_arburst(split111_merge213_arburst[1:0])
    ,.a_arextras(split111_merge213_arextras[(EXTRAS - 1):0])
    ,.a_arid(split111_merge213_arid[(IDWID - 1):0])
    ,.a_arlen(split111_merge213_arlen[7:0])
    ,.a_arready(split111_merge213_arready)
    ,.a_arvalid(split111_merge213_arvalid)
    ,.a_awaddr(split111_merge213_awaddr[31:0])
    ,.a_awburst(split111_merge213_awburst[1:0])
    ,.a_awextras(split111_merge213_awextras[(EXTRAS - 1):0])
    ,.a_awid(split111_merge213_awid[(IDWID - 1):0])
    ,.a_awlen(split111_merge213_awlen[7:0])
    ,.a_awready(split111_merge213_awready)
    ,.a_awvalid(split111_merge213_awvalid)
    ,.a_bid(split111_merge213_bid[(IDWID - 1):0])
    ,.a_bready(split111_merge213_bready)
    ,.a_bresp(split111_merge213_bresp[1:0])
    ,.a_bvalid(split111_merge213_bvalid)
    ,.a_rdata(split111_merge213_rdata[(DWID - 1):0])
    ,.a_rid(split111_merge213_rid[(IDWID - 1):0])
    ,.a_rlast(split111_merge213_rlast)
    ,.a_rready(split111_merge213_rready)
    ,.a_rresp(split111_merge213_rresp[1:0])
    ,.a_rvalid(split111_merge213_rvalid)
    ,.a_wdata(split111_merge213_wdata[(DWID - 1):0])
    ,.a_wlast(split111_merge213_wlast)
    ,.a_wready(split111_merge213_wready)
    ,.a_wstrb(split111_merge213_wstrb[(WSTRB - 1):0])
    ,.a_wvalid(split111_merge213_wvalid)
    ,.b_araddr(split111_merge200_araddr[31:0])
    ,.b_arburst(split111_merge200_arburst[1:0])
    ,.b_arextras(split111_merge200_arextras[(EXTRAS - 1):0])
    ,.b_arid(split111_merge200_arid[(IDWID - 1):0])
    ,.b_arlen(split111_merge200_arlen[7:0])
    ,.b_arready(split111_merge200_arready)
    ,.b_arvalid(split111_merge200_arvalid)
    ,.b_awaddr(split111_merge200_awaddr[31:0])
    ,.b_awburst(split111_merge200_awburst[1:0])
    ,.b_awextras(split111_merge200_awextras[(EXTRAS - 1):0])
    ,.b_awid(split111_merge200_awid[(IDWID - 1):0])
    ,.b_awlen(split111_merge200_awlen[7:0])
    ,.b_awready(split111_merge200_awready)
    ,.b_awvalid(split111_merge200_awvalid)
    ,.b_bid(split111_merge200_bid[(IDWID - 1):0])
    ,.b_bready(split111_merge200_bready)
    ,.b_bresp(split111_merge200_bresp[1:0])
    ,.b_bvalid(split111_merge200_bvalid)
    ,.b_rdata(split111_merge200_rdata[(DWID - 1):0])
    ,.b_rid(split111_merge200_rid[(IDWID - 1):0])
    ,.b_rlast(split111_merge200_rlast)
    ,.b_rready(split111_merge200_rready)
    ,.b_rresp(split111_merge200_rresp[1:0])
    ,.b_rvalid(split111_merge200_rvalid)
    ,.b_wdata(split111_merge200_wdata[(DWID - 1):0])
    ,.b_wlast(split111_merge200_wlast)
    ,.b_wready(split111_merge200_wready)
    ,.b_wstrb(split111_merge200_wstrb[(WSTRB - 1):0])
    ,.b_wvalid(split111_merge200_wvalid)
    ,.c_araddr(split111_merge202_araddr[31:0])
    ,.c_arburst(split111_merge202_arburst[1:0])
    ,.c_arextras(split111_merge202_arextras[(EXTRAS - 1):0])
    ,.c_arid(split111_merge202_arid[(IDWID - 1):0])
    ,.c_arlen(split111_merge202_arlen[7:0])
    ,.c_arready(split111_merge202_arready)
    ,.c_arvalid(split111_merge202_arvalid)
    ,.c_awaddr(split111_merge202_awaddr[31:0])
    ,.c_awburst(split111_merge202_awburst[1:0])
    ,.c_awextras(split111_merge202_awextras[(EXTRAS - 1):0])
    ,.c_awid(split111_merge202_awid[(IDWID - 1):0])
    ,.c_awlen(split111_merge202_awlen[7:0])
    ,.c_awready(split111_merge202_awready)
    ,.c_awvalid(split111_merge202_awvalid)
    ,.c_bid(split111_merge202_bid[(IDWID - 1):0])
    ,.c_bready(split111_merge202_bready)
    ,.c_bresp(split111_merge202_bresp[1:0])
    ,.c_bvalid(split111_merge202_bvalid)
    ,.c_rdata(split111_merge202_rdata[(DWID - 1):0])
    ,.c_rid(split111_merge202_rid[(IDWID - 1):0])
    ,.c_rlast(split111_merge202_rlast)
    ,.c_rready(split111_merge202_rready)
    ,.c_rresp(split111_merge202_rresp[1:0])
    ,.c_rvalid(split111_merge202_rvalid)
    ,.c_wdata(split111_merge202_wdata[(DWID - 1):0])
    ,.c_wlast(split111_merge202_wlast)
    ,.c_wready(split111_merge202_wready)
    ,.c_wstrb(split111_merge202_wstrb[(WSTRB - 1):0])
    ,.c_wvalid(split111_merge202_wvalid)
    ,.d_araddr(split111_merge214_araddr[31:0])
    ,.d_arburst(split111_merge214_arburst[1:0])
    ,.d_arextras(split111_merge214_arextras[(EXTRAS - 1):0])
    ,.d_arid(split111_merge214_arid[(IDWID - 1):0])
    ,.d_arlen(split111_merge214_arlen[7:0])
    ,.d_arready(split111_merge214_arready)
    ,.d_arvalid(split111_merge214_arvalid)
    ,.d_awaddr(split111_merge214_awaddr[31:0])
    ,.d_awburst(split111_merge214_awburst[1:0])
    ,.d_awextras(split111_merge214_awextras[(EXTRAS - 1):0])
    ,.d_awid(split111_merge214_awid[(IDWID - 1):0])
    ,.d_awlen(split111_merge214_awlen[7:0])
    ,.d_awready(split111_merge214_awready)
    ,.d_awvalid(split111_merge214_awvalid)
    ,.d_bid(split111_merge214_bid[(IDWID - 1):0])
    ,.d_bready(split111_merge214_bready)
    ,.d_bresp(split111_merge214_bresp[1:0])
    ,.d_bvalid(split111_merge214_bvalid)
    ,.d_rdata(split111_merge214_rdata[(DWID - 1):0])
    ,.d_rid(split111_merge214_rid[(IDWID - 1):0])
    ,.d_rlast(split111_merge214_rlast)
    ,.d_rready(split111_merge214_rready)
    ,.d_rresp(split111_merge214_rresp[1:0])
    ,.d_rvalid(split111_merge214_rvalid)
    ,.d_wdata(split111_merge214_wdata[(DWID - 1):0])
    ,.d_wlast(split111_merge214_wlast)
    ,.d_wready(split111_merge214_wready)
    ,.d_wstrb(split111_merge214_wstrb[(WSTRB - 1):0])
    ,.d_wvalid(split111_merge214_wvalid)

);

wire [IDWID-1:0] split112_merge215_arid ;
wire [31:0] split112_merge215_araddr ;
wire [7:0] split112_merge215_arlen ;
wire [EXTRAS-1:0] split112_merge215_arextras ;
wire [1:0] split112_merge215_arburst ;
wire split112_merge215_arvalid ;
wire split112_merge215_arready ;
wire [IDWID-1:0] split112_merge215_rid ;
wire [DWID-1:0] split112_merge215_rdata ;
wire [1:0] split112_merge215_rresp ;
wire split112_merge215_rlast ;
wire split112_merge215_rvalid ;
wire split112_merge215_rready ;

wire [IDWID-1:0] split112_merge215_awid ;
wire [31:0] split112_merge215_awaddr ;
wire [7:0] split112_merge215_awlen ;
wire [EXTRAS-1:0] split112_merge215_awextras ;
wire [1:0] split112_merge215_awburst ;
wire split112_merge215_awvalid ;
wire split112_merge215_awready ;
wire [DWID-1:0] split112_merge215_wdata ;
wire [WSTRB-1:0] split112_merge215_wstrb ;
wire split112_merge215_wlast ;
wire split112_merge215_wvalid ;
wire split112_merge215_wready ;
wire [IDWID-1:0] split112_merge215_bid ;
wire [1:0] split112_merge215_bresp ;
wire split112_merge215_bvalid ;
wire split112_merge215_bready ;


wire [IDWID-1:0] split112_merge202_arid ;
wire [31:0] split112_merge202_araddr ;
wire [7:0] split112_merge202_arlen ;
wire [EXTRAS-1:0] split112_merge202_arextras ;
wire [1:0] split112_merge202_arburst ;
wire split112_merge202_arvalid ;
wire split112_merge202_arready ;
wire [IDWID-1:0] split112_merge202_rid ;
wire [DWID-1:0] split112_merge202_rdata ;
wire [1:0] split112_merge202_rresp ;
wire split112_merge202_rlast ;
wire split112_merge202_rvalid ;
wire split112_merge202_rready ;

wire [IDWID-1:0] split112_merge202_awid ;
wire [31:0] split112_merge202_awaddr ;
wire [7:0] split112_merge202_awlen ;
wire [EXTRAS-1:0] split112_merge202_awextras ;
wire [1:0] split112_merge202_awburst ;
wire split112_merge202_awvalid ;
wire split112_merge202_awready ;
wire [DWID-1:0] split112_merge202_wdata ;
wire [WSTRB-1:0] split112_merge202_wstrb ;
wire split112_merge202_wlast ;
wire split112_merge202_wvalid ;
wire split112_merge202_wready ;
wire [IDWID-1:0] split112_merge202_bid ;
wire [1:0] split112_merge202_bresp ;
wire split112_merge202_bvalid ;
wire split112_merge202_bready ;


wire [IDWID-1:0] split112_merge201_arid ;
wire [31:0] split112_merge201_araddr ;
wire [7:0] split112_merge201_arlen ;
wire [EXTRAS-1:0] split112_merge201_arextras ;
wire [1:0] split112_merge201_arburst ;
wire split112_merge201_arvalid ;
wire split112_merge201_arready ;
wire [IDWID-1:0] split112_merge201_rid ;
wire [DWID-1:0] split112_merge201_rdata ;
wire [1:0] split112_merge201_rresp ;
wire split112_merge201_rlast ;
wire split112_merge201_rvalid ;
wire split112_merge201_rready ;

wire [IDWID-1:0] split112_merge201_awid ;
wire [31:0] split112_merge201_awaddr ;
wire [7:0] split112_merge201_awlen ;
wire [EXTRAS-1:0] split112_merge201_awextras ;
wire [1:0] split112_merge201_awburst ;
wire split112_merge201_awvalid ;
wire split112_merge201_awready ;
wire [DWID-1:0] split112_merge201_wdata ;
wire [WSTRB-1:0] split112_merge201_wstrb ;
wire split112_merge201_wlast ;
wire split112_merge201_wvalid ;
wire split112_merge201_wready ;
wire [IDWID-1:0] split112_merge201_bid ;
wire [1:0] split112_merge201_bresp ;
wire split112_merge201_bvalid ;
wire split112_merge201_bready ;


wire [IDWID-1:0] split112_merge210_arid ;
wire [31:0] split112_merge210_araddr ;
wire [7:0] split112_merge210_arlen ;
wire [EXTRAS-1:0] split112_merge210_arextras ;
wire [1:0] split112_merge210_arburst ;
wire split112_merge210_arvalid ;
wire split112_merge210_arready ;
wire [IDWID-1:0] split112_merge210_rid ;
wire [DWID-1:0] split112_merge210_rdata ;
wire [1:0] split112_merge210_rresp ;
wire split112_merge210_rlast ;
wire split112_merge210_rvalid ;
wire split112_merge210_rready ;

wire [IDWID-1:0] split112_merge210_awid ;
wire [31:0] split112_merge210_awaddr ;
wire [7:0] split112_merge210_awlen ;
wire [EXTRAS-1:0] split112_merge210_awextras ;
wire [1:0] split112_merge210_awburst ;
wire split112_merge210_awvalid ;
wire split112_merge210_awready ;
wire [DWID-1:0] split112_merge210_wdata ;
wire [WSTRB-1:0] split112_merge210_wstrb ;
wire split112_merge210_wlast ;
wire split112_merge210_wvalid ;
wire split112_merge210_wready ;
wire [IDWID-1:0] split112_merge210_bid ;
wire [1:0] split112_merge210_bresp ;
wire split112_merge210_bvalid ;
wire split112_merge210_bready ;


axi_4_splitter split112 (
     .clk(clk) ,.rst_n(rst_n)

    ,.araddr(merge12_split112_araddr[31:0])
    ,.arburst(merge12_split112_arburst[1:0])
    ,.arextras(merge12_split112_arextras[(EXTRAS - 1):0])
    ,.arid(merge12_split112_arid[(IDWID - 1):0])
    ,.arlen(merge12_split112_arlen[7:0])
    ,.arready(merge12_split112_arready)
    ,.arvalid(merge12_split112_arvalid)
    ,.awaddr(merge12_split112_awaddr[31:0])
    ,.awburst(merge12_split112_awburst[1:0])
    ,.awextras(merge12_split112_awextras[(EXTRAS - 1):0])
    ,.awid(merge12_split112_awid[3:0])
    ,.awlen(merge12_split112_awlen[7:0])
    ,.awready(merge12_split112_awready)
    ,.awvalid(merge12_split112_awvalid)
    ,.bid(merge12_split112_bid[(IDWID - 1):0])
    ,.bready(merge12_split112_bready)
    ,.bresp(merge12_split112_bresp[1:0])
    ,.bvalid(merge12_split112_bvalid)
    ,.rdata(merge12_split112_rdata[(DWID - 1):0])
    ,.rid(merge12_split112_rid[(IDWID - 1):0])
    ,.rlast(merge12_split112_rlast)
    ,.rready(merge12_split112_rready)
    ,.rresp(merge12_split112_rresp[1:0])
    ,.rvalid(merge12_split112_rvalid)
    ,.wdata(merge12_split112_wdata[(DWID - 1):0])
    ,.wlast(merge12_split112_wlast)
    ,.wready(merge12_split112_wready)
    ,.wstrb(merge12_split112_wstrb[(WSTRB - 1):0])
    ,.wvalid(merge12_split112_wvalid)

    ,.a_araddr(split112_merge215_araddr[31:0])
    ,.a_arburst(split112_merge215_arburst[1:0])
    ,.a_arextras(split112_merge215_arextras[(EXTRAS - 1):0])
    ,.a_arid(split112_merge215_arid[(IDWID - 1):0])
    ,.a_arlen(split112_merge215_arlen[7:0])
    ,.a_arready(split112_merge215_arready)
    ,.a_arvalid(split112_merge215_arvalid)
    ,.a_awaddr(split112_merge215_awaddr[31:0])
    ,.a_awburst(split112_merge215_awburst[1:0])
    ,.a_awextras(split112_merge215_awextras[(EXTRAS - 1):0])
    ,.a_awid(split112_merge215_awid[(IDWID - 1):0])
    ,.a_awlen(split112_merge215_awlen[7:0])
    ,.a_awready(split112_merge215_awready)
    ,.a_awvalid(split112_merge215_awvalid)
    ,.a_bid(split112_merge215_bid[(IDWID - 1):0])
    ,.a_bready(split112_merge215_bready)
    ,.a_bresp(split112_merge215_bresp[1:0])
    ,.a_bvalid(split112_merge215_bvalid)
    ,.a_rdata(split112_merge215_rdata[(DWID - 1):0])
    ,.a_rid(split112_merge215_rid[(IDWID - 1):0])
    ,.a_rlast(split112_merge215_rlast)
    ,.a_rready(split112_merge215_rready)
    ,.a_rresp(split112_merge215_rresp[1:0])
    ,.a_rvalid(split112_merge215_rvalid)
    ,.a_wdata(split112_merge215_wdata[(DWID - 1):0])
    ,.a_wlast(split112_merge215_wlast)
    ,.a_wready(split112_merge215_wready)
    ,.a_wstrb(split112_merge215_wstrb[(WSTRB - 1):0])
    ,.a_wvalid(split112_merge215_wvalid)
    ,.b_araddr(split112_merge202_araddr[31:0])
    ,.b_arburst(split112_merge202_arburst[1:0])
    ,.b_arextras(split112_merge202_arextras[(EXTRAS - 1):0])
    ,.b_arid(split112_merge202_arid[(IDWID - 1):0])
    ,.b_arlen(split112_merge202_arlen[7:0])
    ,.b_arready(split112_merge202_arready)
    ,.b_arvalid(split112_merge202_arvalid)
    ,.b_awaddr(split112_merge202_awaddr[31:0])
    ,.b_awburst(split112_merge202_awburst[1:0])
    ,.b_awextras(split112_merge202_awextras[(EXTRAS - 1):0])
    ,.b_awid(split112_merge202_awid[(IDWID - 1):0])
    ,.b_awlen(split112_merge202_awlen[7:0])
    ,.b_awready(split112_merge202_awready)
    ,.b_awvalid(split112_merge202_awvalid)
    ,.b_bid(split112_merge202_bid[(IDWID - 1):0])
    ,.b_bready(split112_merge202_bready)
    ,.b_bresp(split112_merge202_bresp[1:0])
    ,.b_bvalid(split112_merge202_bvalid)
    ,.b_rdata(split112_merge202_rdata[(DWID - 1):0])
    ,.b_rid(split112_merge202_rid[(IDWID - 1):0])
    ,.b_rlast(split112_merge202_rlast)
    ,.b_rready(split112_merge202_rready)
    ,.b_rresp(split112_merge202_rresp[1:0])
    ,.b_rvalid(split112_merge202_rvalid)
    ,.b_wdata(split112_merge202_wdata[(DWID - 1):0])
    ,.b_wlast(split112_merge202_wlast)
    ,.b_wready(split112_merge202_wready)
    ,.b_wstrb(split112_merge202_wstrb[(WSTRB - 1):0])
    ,.b_wvalid(split112_merge202_wvalid)
    ,.c_araddr(split112_merge201_araddr[31:0])
    ,.c_arburst(split112_merge201_arburst[1:0])
    ,.c_arextras(split112_merge201_arextras[(EXTRAS - 1):0])
    ,.c_arid(split112_merge201_arid[(IDWID - 1):0])
    ,.c_arlen(split112_merge201_arlen[7:0])
    ,.c_arready(split112_merge201_arready)
    ,.c_arvalid(split112_merge201_arvalid)
    ,.c_awaddr(split112_merge201_awaddr[31:0])
    ,.c_awburst(split112_merge201_awburst[1:0])
    ,.c_awextras(split112_merge201_awextras[(EXTRAS - 1):0])
    ,.c_awid(split112_merge201_awid[(IDWID - 1):0])
    ,.c_awlen(split112_merge201_awlen[7:0])
    ,.c_awready(split112_merge201_awready)
    ,.c_awvalid(split112_merge201_awvalid)
    ,.c_bid(split112_merge201_bid[(IDWID - 1):0])
    ,.c_bready(split112_merge201_bready)
    ,.c_bresp(split112_merge201_bresp[1:0])
    ,.c_bvalid(split112_merge201_bvalid)
    ,.c_rdata(split112_merge201_rdata[(DWID - 1):0])
    ,.c_rid(split112_merge201_rid[(IDWID - 1):0])
    ,.c_rlast(split112_merge201_rlast)
    ,.c_rready(split112_merge201_rready)
    ,.c_rresp(split112_merge201_rresp[1:0])
    ,.c_rvalid(split112_merge201_rvalid)
    ,.c_wdata(split112_merge201_wdata[(DWID - 1):0])
    ,.c_wlast(split112_merge201_wlast)
    ,.c_wready(split112_merge201_wready)
    ,.c_wstrb(split112_merge201_wstrb[(WSTRB - 1):0])
    ,.c_wvalid(split112_merge201_wvalid)
    ,.d_araddr(split112_merge210_araddr[31:0])
    ,.d_arburst(split112_merge210_arburst[1:0])
    ,.d_arextras(split112_merge210_arextras[(EXTRAS - 1):0])
    ,.d_arid(split112_merge210_arid[(IDWID - 1):0])
    ,.d_arlen(split112_merge210_arlen[7:0])
    ,.d_arready(split112_merge210_arready)
    ,.d_arvalid(split112_merge210_arvalid)
    ,.d_awaddr(split112_merge210_awaddr[31:0])
    ,.d_awburst(split112_merge210_awburst[1:0])
    ,.d_awextras(split112_merge210_awextras[(EXTRAS - 1):0])
    ,.d_awid(split112_merge210_awid[(IDWID - 1):0])
    ,.d_awlen(split112_merge210_awlen[7:0])
    ,.d_awready(split112_merge210_awready)
    ,.d_awvalid(split112_merge210_awvalid)
    ,.d_bid(split112_merge210_bid[(IDWID - 1):0])
    ,.d_bready(split112_merge210_bready)
    ,.d_bresp(split112_merge210_bresp[1:0])
    ,.d_bvalid(split112_merge210_bvalid)
    ,.d_rdata(split112_merge210_rdata[(DWID - 1):0])
    ,.d_rid(split112_merge210_rid[(IDWID - 1):0])
    ,.d_rlast(split112_merge210_rlast)
    ,.d_rready(split112_merge210_rready)
    ,.d_rresp(split112_merge210_rresp[1:0])
    ,.d_rvalid(split112_merge210_rvalid)
    ,.d_wdata(split112_merge210_wdata[(DWID - 1):0])
    ,.d_wlast(split112_merge210_wlast)
    ,.d_wready(split112_merge210_wready)
    ,.d_wstrb(split112_merge210_wstrb[(WSTRB - 1):0])
    ,.d_wvalid(split112_merge210_wvalid)

);

wire [IDWID-1:0] split113_merge201_arid ;
wire [31:0] split113_merge201_araddr ;
wire [7:0] split113_merge201_arlen ;
wire [EXTRAS-1:0] split113_merge201_arextras ;
wire [1:0] split113_merge201_arburst ;
wire split113_merge201_arvalid ;
wire split113_merge201_arready ;
wire [IDWID-1:0] split113_merge201_rid ;
wire [DWID-1:0] split113_merge201_rdata ;
wire [1:0] split113_merge201_rresp ;
wire split113_merge201_rlast ;
wire split113_merge201_rvalid ;
wire split113_merge201_rready ;

wire [IDWID-1:0] split113_merge201_awid ;
wire [31:0] split113_merge201_awaddr ;
wire [7:0] split113_merge201_awlen ;
wire [EXTRAS-1:0] split113_merge201_awextras ;
wire [1:0] split113_merge201_awburst ;
wire split113_merge201_awvalid ;
wire split113_merge201_awready ;
wire [DWID-1:0] split113_merge201_wdata ;
wire [WSTRB-1:0] split113_merge201_wstrb ;
wire split113_merge201_wlast ;
wire split113_merge201_wvalid ;
wire split113_merge201_wready ;
wire [IDWID-1:0] split113_merge201_bid ;
wire [1:0] split113_merge201_bresp ;
wire split113_merge201_bvalid ;
wire split113_merge201_bready ;


wire [IDWID-1:0] split113_merge206_arid ;
wire [31:0] split113_merge206_araddr ;
wire [7:0] split113_merge206_arlen ;
wire [EXTRAS-1:0] split113_merge206_arextras ;
wire [1:0] split113_merge206_arburst ;
wire split113_merge206_arvalid ;
wire split113_merge206_arready ;
wire [IDWID-1:0] split113_merge206_rid ;
wire [DWID-1:0] split113_merge206_rdata ;
wire [1:0] split113_merge206_rresp ;
wire split113_merge206_rlast ;
wire split113_merge206_rvalid ;
wire split113_merge206_rready ;

wire [IDWID-1:0] split113_merge206_awid ;
wire [31:0] split113_merge206_awaddr ;
wire [7:0] split113_merge206_awlen ;
wire [EXTRAS-1:0] split113_merge206_awextras ;
wire [1:0] split113_merge206_awburst ;
wire split113_merge206_awvalid ;
wire split113_merge206_awready ;
wire [DWID-1:0] split113_merge206_wdata ;
wire [WSTRB-1:0] split113_merge206_wstrb ;
wire split113_merge206_wlast ;
wire split113_merge206_wvalid ;
wire split113_merge206_wready ;
wire [IDWID-1:0] split113_merge206_bid ;
wire [1:0] split113_merge206_bresp ;
wire split113_merge206_bvalid ;
wire split113_merge206_bready ;


wire [IDWID-1:0] split113_merge212_arid ;
wire [31:0] split113_merge212_araddr ;
wire [7:0] split113_merge212_arlen ;
wire [EXTRAS-1:0] split113_merge212_arextras ;
wire [1:0] split113_merge212_arburst ;
wire split113_merge212_arvalid ;
wire split113_merge212_arready ;
wire [IDWID-1:0] split113_merge212_rid ;
wire [DWID-1:0] split113_merge212_rdata ;
wire [1:0] split113_merge212_rresp ;
wire split113_merge212_rlast ;
wire split113_merge212_rvalid ;
wire split113_merge212_rready ;

wire [IDWID-1:0] split113_merge212_awid ;
wire [31:0] split113_merge212_awaddr ;
wire [7:0] split113_merge212_awlen ;
wire [EXTRAS-1:0] split113_merge212_awextras ;
wire [1:0] split113_merge212_awburst ;
wire split113_merge212_awvalid ;
wire split113_merge212_awready ;
wire [DWID-1:0] split113_merge212_wdata ;
wire [WSTRB-1:0] split113_merge212_wstrb ;
wire split113_merge212_wlast ;
wire split113_merge212_wvalid ;
wire split113_merge212_wready ;
wire [IDWID-1:0] split113_merge212_bid ;
wire [1:0] split113_merge212_bresp ;
wire split113_merge212_bvalid ;
wire split113_merge212_bready ;


wire [IDWID-1:0] split113_merge205_arid ;
wire [31:0] split113_merge205_araddr ;
wire [7:0] split113_merge205_arlen ;
wire [EXTRAS-1:0] split113_merge205_arextras ;
wire [1:0] split113_merge205_arburst ;
wire split113_merge205_arvalid ;
wire split113_merge205_arready ;
wire [IDWID-1:0] split113_merge205_rid ;
wire [DWID-1:0] split113_merge205_rdata ;
wire [1:0] split113_merge205_rresp ;
wire split113_merge205_rlast ;
wire split113_merge205_rvalid ;
wire split113_merge205_rready ;

wire [IDWID-1:0] split113_merge205_awid ;
wire [31:0] split113_merge205_awaddr ;
wire [7:0] split113_merge205_awlen ;
wire [EXTRAS-1:0] split113_merge205_awextras ;
wire [1:0] split113_merge205_awburst ;
wire split113_merge205_awvalid ;
wire split113_merge205_awready ;
wire [DWID-1:0] split113_merge205_wdata ;
wire [WSTRB-1:0] split113_merge205_wstrb ;
wire split113_merge205_wlast ;
wire split113_merge205_wvalid ;
wire split113_merge205_wready ;
wire [IDWID-1:0] split113_merge205_bid ;
wire [1:0] split113_merge205_bresp ;
wire split113_merge205_bvalid ;
wire split113_merge205_bready ;


axi_4_splitter split113 (
     .clk(clk) ,.rst_n(rst_n)

    ,.araddr(merge13_split113_araddr[31:0])
    ,.arburst(merge13_split113_arburst[1:0])
    ,.arextras(merge13_split113_arextras[(EXTRAS - 1):0])
    ,.arid(merge13_split113_arid[(IDWID - 1):0])
    ,.arlen(merge13_split113_arlen[7:0])
    ,.arready(merge13_split113_arready)
    ,.arvalid(merge13_split113_arvalid)
    ,.awaddr(merge13_split113_awaddr[31:0])
    ,.awburst(merge13_split113_awburst[1:0])
    ,.awextras(merge13_split113_awextras[(EXTRAS - 1):0])
    ,.awid(merge13_split113_awid[3:0])
    ,.awlen(merge13_split113_awlen[7:0])
    ,.awready(merge13_split113_awready)
    ,.awvalid(merge13_split113_awvalid)
    ,.bid(merge13_split113_bid[(IDWID - 1):0])
    ,.bready(merge13_split113_bready)
    ,.bresp(merge13_split113_bresp[1:0])
    ,.bvalid(merge13_split113_bvalid)
    ,.rdata(merge13_split113_rdata[(DWID - 1):0])
    ,.rid(merge13_split113_rid[(IDWID - 1):0])
    ,.rlast(merge13_split113_rlast)
    ,.rready(merge13_split113_rready)
    ,.rresp(merge13_split113_rresp[1:0])
    ,.rvalid(merge13_split113_rvalid)
    ,.wdata(merge13_split113_wdata[(DWID - 1):0])
    ,.wlast(merge13_split113_wlast)
    ,.wready(merge13_split113_wready)
    ,.wstrb(merge13_split113_wstrb[(WSTRB - 1):0])
    ,.wvalid(merge13_split113_wvalid)

    ,.a_araddr(split113_merge201_araddr[31:0])
    ,.a_arburst(split113_merge201_arburst[1:0])
    ,.a_arextras(split113_merge201_arextras[(EXTRAS - 1):0])
    ,.a_arid(split113_merge201_arid[(IDWID - 1):0])
    ,.a_arlen(split113_merge201_arlen[7:0])
    ,.a_arready(split113_merge201_arready)
    ,.a_arvalid(split113_merge201_arvalid)
    ,.a_awaddr(split113_merge201_awaddr[31:0])
    ,.a_awburst(split113_merge201_awburst[1:0])
    ,.a_awextras(split113_merge201_awextras[(EXTRAS - 1):0])
    ,.a_awid(split113_merge201_awid[(IDWID - 1):0])
    ,.a_awlen(split113_merge201_awlen[7:0])
    ,.a_awready(split113_merge201_awready)
    ,.a_awvalid(split113_merge201_awvalid)
    ,.a_bid(split113_merge201_bid[(IDWID - 1):0])
    ,.a_bready(split113_merge201_bready)
    ,.a_bresp(split113_merge201_bresp[1:0])
    ,.a_bvalid(split113_merge201_bvalid)
    ,.a_rdata(split113_merge201_rdata[(DWID - 1):0])
    ,.a_rid(split113_merge201_rid[(IDWID - 1):0])
    ,.a_rlast(split113_merge201_rlast)
    ,.a_rready(split113_merge201_rready)
    ,.a_rresp(split113_merge201_rresp[1:0])
    ,.a_rvalid(split113_merge201_rvalid)
    ,.a_wdata(split113_merge201_wdata[(DWID - 1):0])
    ,.a_wlast(split113_merge201_wlast)
    ,.a_wready(split113_merge201_wready)
    ,.a_wstrb(split113_merge201_wstrb[(WSTRB - 1):0])
    ,.a_wvalid(split113_merge201_wvalid)
    ,.b_araddr(split113_merge206_araddr[31:0])
    ,.b_arburst(split113_merge206_arburst[1:0])
    ,.b_arextras(split113_merge206_arextras[(EXTRAS - 1):0])
    ,.b_arid(split113_merge206_arid[(IDWID - 1):0])
    ,.b_arlen(split113_merge206_arlen[7:0])
    ,.b_arready(split113_merge206_arready)
    ,.b_arvalid(split113_merge206_arvalid)
    ,.b_awaddr(split113_merge206_awaddr[31:0])
    ,.b_awburst(split113_merge206_awburst[1:0])
    ,.b_awextras(split113_merge206_awextras[(EXTRAS - 1):0])
    ,.b_awid(split113_merge206_awid[(IDWID - 1):0])
    ,.b_awlen(split113_merge206_awlen[7:0])
    ,.b_awready(split113_merge206_awready)
    ,.b_awvalid(split113_merge206_awvalid)
    ,.b_bid(split113_merge206_bid[(IDWID - 1):0])
    ,.b_bready(split113_merge206_bready)
    ,.b_bresp(split113_merge206_bresp[1:0])
    ,.b_bvalid(split113_merge206_bvalid)
    ,.b_rdata(split113_merge206_rdata[(DWID - 1):0])
    ,.b_rid(split113_merge206_rid[(IDWID - 1):0])
    ,.b_rlast(split113_merge206_rlast)
    ,.b_rready(split113_merge206_rready)
    ,.b_rresp(split113_merge206_rresp[1:0])
    ,.b_rvalid(split113_merge206_rvalid)
    ,.b_wdata(split113_merge206_wdata[(DWID - 1):0])
    ,.b_wlast(split113_merge206_wlast)
    ,.b_wready(split113_merge206_wready)
    ,.b_wstrb(split113_merge206_wstrb[(WSTRB - 1):0])
    ,.b_wvalid(split113_merge206_wvalid)
    ,.c_araddr(split113_merge212_araddr[31:0])
    ,.c_arburst(split113_merge212_arburst[1:0])
    ,.c_arextras(split113_merge212_arextras[(EXTRAS - 1):0])
    ,.c_arid(split113_merge212_arid[(IDWID - 1):0])
    ,.c_arlen(split113_merge212_arlen[7:0])
    ,.c_arready(split113_merge212_arready)
    ,.c_arvalid(split113_merge212_arvalid)
    ,.c_awaddr(split113_merge212_awaddr[31:0])
    ,.c_awburst(split113_merge212_awburst[1:0])
    ,.c_awextras(split113_merge212_awextras[(EXTRAS - 1):0])
    ,.c_awid(split113_merge212_awid[(IDWID - 1):0])
    ,.c_awlen(split113_merge212_awlen[7:0])
    ,.c_awready(split113_merge212_awready)
    ,.c_awvalid(split113_merge212_awvalid)
    ,.c_bid(split113_merge212_bid[(IDWID - 1):0])
    ,.c_bready(split113_merge212_bready)
    ,.c_bresp(split113_merge212_bresp[1:0])
    ,.c_bvalid(split113_merge212_bvalid)
    ,.c_rdata(split113_merge212_rdata[(DWID - 1):0])
    ,.c_rid(split113_merge212_rid[(IDWID - 1):0])
    ,.c_rlast(split113_merge212_rlast)
    ,.c_rready(split113_merge212_rready)
    ,.c_rresp(split113_merge212_rresp[1:0])
    ,.c_rvalid(split113_merge212_rvalid)
    ,.c_wdata(split113_merge212_wdata[(DWID - 1):0])
    ,.c_wlast(split113_merge212_wlast)
    ,.c_wready(split113_merge212_wready)
    ,.c_wstrb(split113_merge212_wstrb[(WSTRB - 1):0])
    ,.c_wvalid(split113_merge212_wvalid)
    ,.d_araddr(split113_merge205_araddr[31:0])
    ,.d_arburst(split113_merge205_arburst[1:0])
    ,.d_arextras(split113_merge205_arextras[(EXTRAS - 1):0])
    ,.d_arid(split113_merge205_arid[(IDWID - 1):0])
    ,.d_arlen(split113_merge205_arlen[7:0])
    ,.d_arready(split113_merge205_arready)
    ,.d_arvalid(split113_merge205_arvalid)
    ,.d_awaddr(split113_merge205_awaddr[31:0])
    ,.d_awburst(split113_merge205_awburst[1:0])
    ,.d_awextras(split113_merge205_awextras[(EXTRAS - 1):0])
    ,.d_awid(split113_merge205_awid[(IDWID - 1):0])
    ,.d_awlen(split113_merge205_awlen[7:0])
    ,.d_awready(split113_merge205_awready)
    ,.d_awvalid(split113_merge205_awvalid)
    ,.d_bid(split113_merge205_bid[(IDWID - 1):0])
    ,.d_bready(split113_merge205_bready)
    ,.d_bresp(split113_merge205_bresp[1:0])
    ,.d_bvalid(split113_merge205_bvalid)
    ,.d_rdata(split113_merge205_rdata[(DWID - 1):0])
    ,.d_rid(split113_merge205_rid[(IDWID - 1):0])
    ,.d_rlast(split113_merge205_rlast)
    ,.d_rready(split113_merge205_rready)
    ,.d_rresp(split113_merge205_rresp[1:0])
    ,.d_rvalid(split113_merge205_rvalid)
    ,.d_wdata(split113_merge205_wdata[(DWID - 1):0])
    ,.d_wlast(split113_merge205_wlast)
    ,.d_wready(split113_merge205_wready)
    ,.d_wstrb(split113_merge205_wstrb[(WSTRB - 1):0])
    ,.d_wvalid(split113_merge205_wvalid)

);

wire [IDWID-1:0] split114_merge208_arid ;
wire [31:0] split114_merge208_araddr ;
wire [7:0] split114_merge208_arlen ;
wire [EXTRAS-1:0] split114_merge208_arextras ;
wire [1:0] split114_merge208_arburst ;
wire split114_merge208_arvalid ;
wire split114_merge208_arready ;
wire [IDWID-1:0] split114_merge208_rid ;
wire [DWID-1:0] split114_merge208_rdata ;
wire [1:0] split114_merge208_rresp ;
wire split114_merge208_rlast ;
wire split114_merge208_rvalid ;
wire split114_merge208_rready ;

wire [IDWID-1:0] split114_merge208_awid ;
wire [31:0] split114_merge208_awaddr ;
wire [7:0] split114_merge208_awlen ;
wire [EXTRAS-1:0] split114_merge208_awextras ;
wire [1:0] split114_merge208_awburst ;
wire split114_merge208_awvalid ;
wire split114_merge208_awready ;
wire [DWID-1:0] split114_merge208_wdata ;
wire [WSTRB-1:0] split114_merge208_wstrb ;
wire split114_merge208_wlast ;
wire split114_merge208_wvalid ;
wire split114_merge208_wready ;
wire [IDWID-1:0] split114_merge208_bid ;
wire [1:0] split114_merge208_bresp ;
wire split114_merge208_bvalid ;
wire split114_merge208_bready ;


wire [IDWID-1:0] split114_merge210_arid ;
wire [31:0] split114_merge210_araddr ;
wire [7:0] split114_merge210_arlen ;
wire [EXTRAS-1:0] split114_merge210_arextras ;
wire [1:0] split114_merge210_arburst ;
wire split114_merge210_arvalid ;
wire split114_merge210_arready ;
wire [IDWID-1:0] split114_merge210_rid ;
wire [DWID-1:0] split114_merge210_rdata ;
wire [1:0] split114_merge210_rresp ;
wire split114_merge210_rlast ;
wire split114_merge210_rvalid ;
wire split114_merge210_rready ;

wire [IDWID-1:0] split114_merge210_awid ;
wire [31:0] split114_merge210_awaddr ;
wire [7:0] split114_merge210_awlen ;
wire [EXTRAS-1:0] split114_merge210_awextras ;
wire [1:0] split114_merge210_awburst ;
wire split114_merge210_awvalid ;
wire split114_merge210_awready ;
wire [DWID-1:0] split114_merge210_wdata ;
wire [WSTRB-1:0] split114_merge210_wstrb ;
wire split114_merge210_wlast ;
wire split114_merge210_wvalid ;
wire split114_merge210_wready ;
wire [IDWID-1:0] split114_merge210_bid ;
wire [1:0] split114_merge210_bresp ;
wire split114_merge210_bvalid ;
wire split114_merge210_bready ;


wire [IDWID-1:0] split114_merge215_arid ;
wire [31:0] split114_merge215_araddr ;
wire [7:0] split114_merge215_arlen ;
wire [EXTRAS-1:0] split114_merge215_arextras ;
wire [1:0] split114_merge215_arburst ;
wire split114_merge215_arvalid ;
wire split114_merge215_arready ;
wire [IDWID-1:0] split114_merge215_rid ;
wire [DWID-1:0] split114_merge215_rdata ;
wire [1:0] split114_merge215_rresp ;
wire split114_merge215_rlast ;
wire split114_merge215_rvalid ;
wire split114_merge215_rready ;

wire [IDWID-1:0] split114_merge215_awid ;
wire [31:0] split114_merge215_awaddr ;
wire [7:0] split114_merge215_awlen ;
wire [EXTRAS-1:0] split114_merge215_awextras ;
wire [1:0] split114_merge215_awburst ;
wire split114_merge215_awvalid ;
wire split114_merge215_awready ;
wire [DWID-1:0] split114_merge215_wdata ;
wire [WSTRB-1:0] split114_merge215_wstrb ;
wire split114_merge215_wlast ;
wire split114_merge215_wvalid ;
wire split114_merge215_wready ;
wire [IDWID-1:0] split114_merge215_bid ;
wire [1:0] split114_merge215_bresp ;
wire split114_merge215_bvalid ;
wire split114_merge215_bready ;


wire [IDWID-1:0] split114_merge204_arid ;
wire [31:0] split114_merge204_araddr ;
wire [7:0] split114_merge204_arlen ;
wire [EXTRAS-1:0] split114_merge204_arextras ;
wire [1:0] split114_merge204_arburst ;
wire split114_merge204_arvalid ;
wire split114_merge204_arready ;
wire [IDWID-1:0] split114_merge204_rid ;
wire [DWID-1:0] split114_merge204_rdata ;
wire [1:0] split114_merge204_rresp ;
wire split114_merge204_rlast ;
wire split114_merge204_rvalid ;
wire split114_merge204_rready ;

wire [IDWID-1:0] split114_merge204_awid ;
wire [31:0] split114_merge204_awaddr ;
wire [7:0] split114_merge204_awlen ;
wire [EXTRAS-1:0] split114_merge204_awextras ;
wire [1:0] split114_merge204_awburst ;
wire split114_merge204_awvalid ;
wire split114_merge204_awready ;
wire [DWID-1:0] split114_merge204_wdata ;
wire [WSTRB-1:0] split114_merge204_wstrb ;
wire split114_merge204_wlast ;
wire split114_merge204_wvalid ;
wire split114_merge204_wready ;
wire [IDWID-1:0] split114_merge204_bid ;
wire [1:0] split114_merge204_bresp ;
wire split114_merge204_bvalid ;
wire split114_merge204_bready ;


axi_4_splitter split114 (
     .clk(clk) ,.rst_n(rst_n)

    ,.araddr(merge14_split114_araddr[31:0])
    ,.arburst(merge14_split114_arburst[1:0])
    ,.arextras(merge14_split114_arextras[(EXTRAS - 1):0])
    ,.arid(merge14_split114_arid[(IDWID - 1):0])
    ,.arlen(merge14_split114_arlen[7:0])
    ,.arready(merge14_split114_arready)
    ,.arvalid(merge14_split114_arvalid)
    ,.awaddr(merge14_split114_awaddr[31:0])
    ,.awburst(merge14_split114_awburst[1:0])
    ,.awextras(merge14_split114_awextras[(EXTRAS - 1):0])
    ,.awid(merge14_split114_awid[3:0])
    ,.awlen(merge14_split114_awlen[7:0])
    ,.awready(merge14_split114_awready)
    ,.awvalid(merge14_split114_awvalid)
    ,.bid(merge14_split114_bid[(IDWID - 1):0])
    ,.bready(merge14_split114_bready)
    ,.bresp(merge14_split114_bresp[1:0])
    ,.bvalid(merge14_split114_bvalid)
    ,.rdata(merge14_split114_rdata[(DWID - 1):0])
    ,.rid(merge14_split114_rid[(IDWID - 1):0])
    ,.rlast(merge14_split114_rlast)
    ,.rready(merge14_split114_rready)
    ,.rresp(merge14_split114_rresp[1:0])
    ,.rvalid(merge14_split114_rvalid)
    ,.wdata(merge14_split114_wdata[(DWID - 1):0])
    ,.wlast(merge14_split114_wlast)
    ,.wready(merge14_split114_wready)
    ,.wstrb(merge14_split114_wstrb[(WSTRB - 1):0])
    ,.wvalid(merge14_split114_wvalid)

    ,.a_araddr(split114_merge208_araddr[31:0])
    ,.a_arburst(split114_merge208_arburst[1:0])
    ,.a_arextras(split114_merge208_arextras[(EXTRAS - 1):0])
    ,.a_arid(split114_merge208_arid[(IDWID - 1):0])
    ,.a_arlen(split114_merge208_arlen[7:0])
    ,.a_arready(split114_merge208_arready)
    ,.a_arvalid(split114_merge208_arvalid)
    ,.a_awaddr(split114_merge208_awaddr[31:0])
    ,.a_awburst(split114_merge208_awburst[1:0])
    ,.a_awextras(split114_merge208_awextras[(EXTRAS - 1):0])
    ,.a_awid(split114_merge208_awid[(IDWID - 1):0])
    ,.a_awlen(split114_merge208_awlen[7:0])
    ,.a_awready(split114_merge208_awready)
    ,.a_awvalid(split114_merge208_awvalid)
    ,.a_bid(split114_merge208_bid[(IDWID - 1):0])
    ,.a_bready(split114_merge208_bready)
    ,.a_bresp(split114_merge208_bresp[1:0])
    ,.a_bvalid(split114_merge208_bvalid)
    ,.a_rdata(split114_merge208_rdata[(DWID - 1):0])
    ,.a_rid(split114_merge208_rid[(IDWID - 1):0])
    ,.a_rlast(split114_merge208_rlast)
    ,.a_rready(split114_merge208_rready)
    ,.a_rresp(split114_merge208_rresp[1:0])
    ,.a_rvalid(split114_merge208_rvalid)
    ,.a_wdata(split114_merge208_wdata[(DWID - 1):0])
    ,.a_wlast(split114_merge208_wlast)
    ,.a_wready(split114_merge208_wready)
    ,.a_wstrb(split114_merge208_wstrb[(WSTRB - 1):0])
    ,.a_wvalid(split114_merge208_wvalid)
    ,.b_araddr(split114_merge210_araddr[31:0])
    ,.b_arburst(split114_merge210_arburst[1:0])
    ,.b_arextras(split114_merge210_arextras[(EXTRAS - 1):0])
    ,.b_arid(split114_merge210_arid[(IDWID - 1):0])
    ,.b_arlen(split114_merge210_arlen[7:0])
    ,.b_arready(split114_merge210_arready)
    ,.b_arvalid(split114_merge210_arvalid)
    ,.b_awaddr(split114_merge210_awaddr[31:0])
    ,.b_awburst(split114_merge210_awburst[1:0])
    ,.b_awextras(split114_merge210_awextras[(EXTRAS - 1):0])
    ,.b_awid(split114_merge210_awid[(IDWID - 1):0])
    ,.b_awlen(split114_merge210_awlen[7:0])
    ,.b_awready(split114_merge210_awready)
    ,.b_awvalid(split114_merge210_awvalid)
    ,.b_bid(split114_merge210_bid[(IDWID - 1):0])
    ,.b_bready(split114_merge210_bready)
    ,.b_bresp(split114_merge210_bresp[1:0])
    ,.b_bvalid(split114_merge210_bvalid)
    ,.b_rdata(split114_merge210_rdata[(DWID - 1):0])
    ,.b_rid(split114_merge210_rid[(IDWID - 1):0])
    ,.b_rlast(split114_merge210_rlast)
    ,.b_rready(split114_merge210_rready)
    ,.b_rresp(split114_merge210_rresp[1:0])
    ,.b_rvalid(split114_merge210_rvalid)
    ,.b_wdata(split114_merge210_wdata[(DWID - 1):0])
    ,.b_wlast(split114_merge210_wlast)
    ,.b_wready(split114_merge210_wready)
    ,.b_wstrb(split114_merge210_wstrb[(WSTRB - 1):0])
    ,.b_wvalid(split114_merge210_wvalid)
    ,.c_araddr(split114_merge215_araddr[31:0])
    ,.c_arburst(split114_merge215_arburst[1:0])
    ,.c_arextras(split114_merge215_arextras[(EXTRAS - 1):0])
    ,.c_arid(split114_merge215_arid[(IDWID - 1):0])
    ,.c_arlen(split114_merge215_arlen[7:0])
    ,.c_arready(split114_merge215_arready)
    ,.c_arvalid(split114_merge215_arvalid)
    ,.c_awaddr(split114_merge215_awaddr[31:0])
    ,.c_awburst(split114_merge215_awburst[1:0])
    ,.c_awextras(split114_merge215_awextras[(EXTRAS - 1):0])
    ,.c_awid(split114_merge215_awid[(IDWID - 1):0])
    ,.c_awlen(split114_merge215_awlen[7:0])
    ,.c_awready(split114_merge215_awready)
    ,.c_awvalid(split114_merge215_awvalid)
    ,.c_bid(split114_merge215_bid[(IDWID - 1):0])
    ,.c_bready(split114_merge215_bready)
    ,.c_bresp(split114_merge215_bresp[1:0])
    ,.c_bvalid(split114_merge215_bvalid)
    ,.c_rdata(split114_merge215_rdata[(DWID - 1):0])
    ,.c_rid(split114_merge215_rid[(IDWID - 1):0])
    ,.c_rlast(split114_merge215_rlast)
    ,.c_rready(split114_merge215_rready)
    ,.c_rresp(split114_merge215_rresp[1:0])
    ,.c_rvalid(split114_merge215_rvalid)
    ,.c_wdata(split114_merge215_wdata[(DWID - 1):0])
    ,.c_wlast(split114_merge215_wlast)
    ,.c_wready(split114_merge215_wready)
    ,.c_wstrb(split114_merge215_wstrb[(WSTRB - 1):0])
    ,.c_wvalid(split114_merge215_wvalid)
    ,.d_araddr(split114_merge204_araddr[31:0])
    ,.d_arburst(split114_merge204_arburst[1:0])
    ,.d_arextras(split114_merge204_arextras[(EXTRAS - 1):0])
    ,.d_arid(split114_merge204_arid[(IDWID - 1):0])
    ,.d_arlen(split114_merge204_arlen[7:0])
    ,.d_arready(split114_merge204_arready)
    ,.d_arvalid(split114_merge204_arvalid)
    ,.d_awaddr(split114_merge204_awaddr[31:0])
    ,.d_awburst(split114_merge204_awburst[1:0])
    ,.d_awextras(split114_merge204_awextras[(EXTRAS - 1):0])
    ,.d_awid(split114_merge204_awid[(IDWID - 1):0])
    ,.d_awlen(split114_merge204_awlen[7:0])
    ,.d_awready(split114_merge204_awready)
    ,.d_awvalid(split114_merge204_awvalid)
    ,.d_bid(split114_merge204_bid[(IDWID - 1):0])
    ,.d_bready(split114_merge204_bready)
    ,.d_bresp(split114_merge204_bresp[1:0])
    ,.d_bvalid(split114_merge204_bvalid)
    ,.d_rdata(split114_merge204_rdata[(DWID - 1):0])
    ,.d_rid(split114_merge204_rid[(IDWID - 1):0])
    ,.d_rlast(split114_merge204_rlast)
    ,.d_rready(split114_merge204_rready)
    ,.d_rresp(split114_merge204_rresp[1:0])
    ,.d_rvalid(split114_merge204_rvalid)
    ,.d_wdata(split114_merge204_wdata[(DWID - 1):0])
    ,.d_wlast(split114_merge204_wlast)
    ,.d_wready(split114_merge204_wready)
    ,.d_wstrb(split114_merge204_wstrb[(WSTRB - 1):0])
    ,.d_wvalid(split114_merge204_wvalid)

);

wire [IDWID-1:0] split115_merge210_arid ;
wire [31:0] split115_merge210_araddr ;
wire [7:0] split115_merge210_arlen ;
wire [EXTRAS-1:0] split115_merge210_arextras ;
wire [1:0] split115_merge210_arburst ;
wire split115_merge210_arvalid ;
wire split115_merge210_arready ;
wire [IDWID-1:0] split115_merge210_rid ;
wire [DWID-1:0] split115_merge210_rdata ;
wire [1:0] split115_merge210_rresp ;
wire split115_merge210_rlast ;
wire split115_merge210_rvalid ;
wire split115_merge210_rready ;

wire [IDWID-1:0] split115_merge210_awid ;
wire [31:0] split115_merge210_awaddr ;
wire [7:0] split115_merge210_awlen ;
wire [EXTRAS-1:0] split115_merge210_awextras ;
wire [1:0] split115_merge210_awburst ;
wire split115_merge210_awvalid ;
wire split115_merge210_awready ;
wire [DWID-1:0] split115_merge210_wdata ;
wire [WSTRB-1:0] split115_merge210_wstrb ;
wire split115_merge210_wlast ;
wire split115_merge210_wvalid ;
wire split115_merge210_wready ;
wire [IDWID-1:0] split115_merge210_bid ;
wire [1:0] split115_merge210_bresp ;
wire split115_merge210_bvalid ;
wire split115_merge210_bready ;


wire [IDWID-1:0] split115_merge207_arid ;
wire [31:0] split115_merge207_araddr ;
wire [7:0] split115_merge207_arlen ;
wire [EXTRAS-1:0] split115_merge207_arextras ;
wire [1:0] split115_merge207_arburst ;
wire split115_merge207_arvalid ;
wire split115_merge207_arready ;
wire [IDWID-1:0] split115_merge207_rid ;
wire [DWID-1:0] split115_merge207_rdata ;
wire [1:0] split115_merge207_rresp ;
wire split115_merge207_rlast ;
wire split115_merge207_rvalid ;
wire split115_merge207_rready ;

wire [IDWID-1:0] split115_merge207_awid ;
wire [31:0] split115_merge207_awaddr ;
wire [7:0] split115_merge207_awlen ;
wire [EXTRAS-1:0] split115_merge207_awextras ;
wire [1:0] split115_merge207_awburst ;
wire split115_merge207_awvalid ;
wire split115_merge207_awready ;
wire [DWID-1:0] split115_merge207_wdata ;
wire [WSTRB-1:0] split115_merge207_wstrb ;
wire split115_merge207_wlast ;
wire split115_merge207_wvalid ;
wire split115_merge207_wready ;
wire [IDWID-1:0] split115_merge207_bid ;
wire [1:0] split115_merge207_bresp ;
wire split115_merge207_bvalid ;
wire split115_merge207_bready ;


wire [IDWID-1:0] split115_merge214_arid ;
wire [31:0] split115_merge214_araddr ;
wire [7:0] split115_merge214_arlen ;
wire [EXTRAS-1:0] split115_merge214_arextras ;
wire [1:0] split115_merge214_arburst ;
wire split115_merge214_arvalid ;
wire split115_merge214_arready ;
wire [IDWID-1:0] split115_merge214_rid ;
wire [DWID-1:0] split115_merge214_rdata ;
wire [1:0] split115_merge214_rresp ;
wire split115_merge214_rlast ;
wire split115_merge214_rvalid ;
wire split115_merge214_rready ;

wire [IDWID-1:0] split115_merge214_awid ;
wire [31:0] split115_merge214_awaddr ;
wire [7:0] split115_merge214_awlen ;
wire [EXTRAS-1:0] split115_merge214_awextras ;
wire [1:0] split115_merge214_awburst ;
wire split115_merge214_awvalid ;
wire split115_merge214_awready ;
wire [DWID-1:0] split115_merge214_wdata ;
wire [WSTRB-1:0] split115_merge214_wstrb ;
wire split115_merge214_wlast ;
wire split115_merge214_wvalid ;
wire split115_merge214_wready ;
wire [IDWID-1:0] split115_merge214_bid ;
wire [1:0] split115_merge214_bresp ;
wire split115_merge214_bvalid ;
wire split115_merge214_bready ;


wire [IDWID-1:0] split115_merge208_arid ;
wire [31:0] split115_merge208_araddr ;
wire [7:0] split115_merge208_arlen ;
wire [EXTRAS-1:0] split115_merge208_arextras ;
wire [1:0] split115_merge208_arburst ;
wire split115_merge208_arvalid ;
wire split115_merge208_arready ;
wire [IDWID-1:0] split115_merge208_rid ;
wire [DWID-1:0] split115_merge208_rdata ;
wire [1:0] split115_merge208_rresp ;
wire split115_merge208_rlast ;
wire split115_merge208_rvalid ;
wire split115_merge208_rready ;

wire [IDWID-1:0] split115_merge208_awid ;
wire [31:0] split115_merge208_awaddr ;
wire [7:0] split115_merge208_awlen ;
wire [EXTRAS-1:0] split115_merge208_awextras ;
wire [1:0] split115_merge208_awburst ;
wire split115_merge208_awvalid ;
wire split115_merge208_awready ;
wire [DWID-1:0] split115_merge208_wdata ;
wire [WSTRB-1:0] split115_merge208_wstrb ;
wire split115_merge208_wlast ;
wire split115_merge208_wvalid ;
wire split115_merge208_wready ;
wire [IDWID-1:0] split115_merge208_bid ;
wire [1:0] split115_merge208_bresp ;
wire split115_merge208_bvalid ;
wire split115_merge208_bready ;


axi_4_splitter split115 (
     .clk(clk) ,.rst_n(rst_n)

    ,.araddr(merge15_split115_araddr[31:0])
    ,.arburst(merge15_split115_arburst[1:0])
    ,.arextras(merge15_split115_arextras[(EXTRAS - 1):0])
    ,.arid(merge15_split115_arid[(IDWID - 1):0])
    ,.arlen(merge15_split115_arlen[7:0])
    ,.arready(merge15_split115_arready)
    ,.arvalid(merge15_split115_arvalid)
    ,.awaddr(merge15_split115_awaddr[31:0])
    ,.awburst(merge15_split115_awburst[1:0])
    ,.awextras(merge15_split115_awextras[(EXTRAS - 1):0])
    ,.awid(merge15_split115_awid[3:0])
    ,.awlen(merge15_split115_awlen[7:0])
    ,.awready(merge15_split115_awready)
    ,.awvalid(merge15_split115_awvalid)
    ,.bid(merge15_split115_bid[(IDWID - 1):0])
    ,.bready(merge15_split115_bready)
    ,.bresp(merge15_split115_bresp[1:0])
    ,.bvalid(merge15_split115_bvalid)
    ,.rdata(merge15_split115_rdata[(DWID - 1):0])
    ,.rid(merge15_split115_rid[(IDWID - 1):0])
    ,.rlast(merge15_split115_rlast)
    ,.rready(merge15_split115_rready)
    ,.rresp(merge15_split115_rresp[1:0])
    ,.rvalid(merge15_split115_rvalid)
    ,.wdata(merge15_split115_wdata[(DWID - 1):0])
    ,.wlast(merge15_split115_wlast)
    ,.wready(merge15_split115_wready)
    ,.wstrb(merge15_split115_wstrb[(WSTRB - 1):0])
    ,.wvalid(merge15_split115_wvalid)

    ,.a_araddr(split115_merge210_araddr[31:0])
    ,.a_arburst(split115_merge210_arburst[1:0])
    ,.a_arextras(split115_merge210_arextras[(EXTRAS - 1):0])
    ,.a_arid(split115_merge210_arid[(IDWID - 1):0])
    ,.a_arlen(split115_merge210_arlen[7:0])
    ,.a_arready(split115_merge210_arready)
    ,.a_arvalid(split115_merge210_arvalid)
    ,.a_awaddr(split115_merge210_awaddr[31:0])
    ,.a_awburst(split115_merge210_awburst[1:0])
    ,.a_awextras(split115_merge210_awextras[(EXTRAS - 1):0])
    ,.a_awid(split115_merge210_awid[(IDWID - 1):0])
    ,.a_awlen(split115_merge210_awlen[7:0])
    ,.a_awready(split115_merge210_awready)
    ,.a_awvalid(split115_merge210_awvalid)
    ,.a_bid(split115_merge210_bid[(IDWID - 1):0])
    ,.a_bready(split115_merge210_bready)
    ,.a_bresp(split115_merge210_bresp[1:0])
    ,.a_bvalid(split115_merge210_bvalid)
    ,.a_rdata(split115_merge210_rdata[(DWID - 1):0])
    ,.a_rid(split115_merge210_rid[(IDWID - 1):0])
    ,.a_rlast(split115_merge210_rlast)
    ,.a_rready(split115_merge210_rready)
    ,.a_rresp(split115_merge210_rresp[1:0])
    ,.a_rvalid(split115_merge210_rvalid)
    ,.a_wdata(split115_merge210_wdata[(DWID - 1):0])
    ,.a_wlast(split115_merge210_wlast)
    ,.a_wready(split115_merge210_wready)
    ,.a_wstrb(split115_merge210_wstrb[(WSTRB - 1):0])
    ,.a_wvalid(split115_merge210_wvalid)
    ,.b_araddr(split115_merge207_araddr[31:0])
    ,.b_arburst(split115_merge207_arburst[1:0])
    ,.b_arextras(split115_merge207_arextras[(EXTRAS - 1):0])
    ,.b_arid(split115_merge207_arid[(IDWID - 1):0])
    ,.b_arlen(split115_merge207_arlen[7:0])
    ,.b_arready(split115_merge207_arready)
    ,.b_arvalid(split115_merge207_arvalid)
    ,.b_awaddr(split115_merge207_awaddr[31:0])
    ,.b_awburst(split115_merge207_awburst[1:0])
    ,.b_awextras(split115_merge207_awextras[(EXTRAS - 1):0])
    ,.b_awid(split115_merge207_awid[(IDWID - 1):0])
    ,.b_awlen(split115_merge207_awlen[7:0])
    ,.b_awready(split115_merge207_awready)
    ,.b_awvalid(split115_merge207_awvalid)
    ,.b_bid(split115_merge207_bid[(IDWID - 1):0])
    ,.b_bready(split115_merge207_bready)
    ,.b_bresp(split115_merge207_bresp[1:0])
    ,.b_bvalid(split115_merge207_bvalid)
    ,.b_rdata(split115_merge207_rdata[(DWID - 1):0])
    ,.b_rid(split115_merge207_rid[(IDWID - 1):0])
    ,.b_rlast(split115_merge207_rlast)
    ,.b_rready(split115_merge207_rready)
    ,.b_rresp(split115_merge207_rresp[1:0])
    ,.b_rvalid(split115_merge207_rvalid)
    ,.b_wdata(split115_merge207_wdata[(DWID - 1):0])
    ,.b_wlast(split115_merge207_wlast)
    ,.b_wready(split115_merge207_wready)
    ,.b_wstrb(split115_merge207_wstrb[(WSTRB - 1):0])
    ,.b_wvalid(split115_merge207_wvalid)
    ,.c_araddr(split115_merge214_araddr[31:0])
    ,.c_arburst(split115_merge214_arburst[1:0])
    ,.c_arextras(split115_merge214_arextras[(EXTRAS - 1):0])
    ,.c_arid(split115_merge214_arid[(IDWID - 1):0])
    ,.c_arlen(split115_merge214_arlen[7:0])
    ,.c_arready(split115_merge214_arready)
    ,.c_arvalid(split115_merge214_arvalid)
    ,.c_awaddr(split115_merge214_awaddr[31:0])
    ,.c_awburst(split115_merge214_awburst[1:0])
    ,.c_awextras(split115_merge214_awextras[(EXTRAS - 1):0])
    ,.c_awid(split115_merge214_awid[(IDWID - 1):0])
    ,.c_awlen(split115_merge214_awlen[7:0])
    ,.c_awready(split115_merge214_awready)
    ,.c_awvalid(split115_merge214_awvalid)
    ,.c_bid(split115_merge214_bid[(IDWID - 1):0])
    ,.c_bready(split115_merge214_bready)
    ,.c_bresp(split115_merge214_bresp[1:0])
    ,.c_bvalid(split115_merge214_bvalid)
    ,.c_rdata(split115_merge214_rdata[(DWID - 1):0])
    ,.c_rid(split115_merge214_rid[(IDWID - 1):0])
    ,.c_rlast(split115_merge214_rlast)
    ,.c_rready(split115_merge214_rready)
    ,.c_rresp(split115_merge214_rresp[1:0])
    ,.c_rvalid(split115_merge214_rvalid)
    ,.c_wdata(split115_merge214_wdata[(DWID - 1):0])
    ,.c_wlast(split115_merge214_wlast)
    ,.c_wready(split115_merge214_wready)
    ,.c_wstrb(split115_merge214_wstrb[(WSTRB - 1):0])
    ,.c_wvalid(split115_merge214_wvalid)
    ,.d_araddr(split115_merge208_araddr[31:0])
    ,.d_arburst(split115_merge208_arburst[1:0])
    ,.d_arextras(split115_merge208_arextras[(EXTRAS - 1):0])
    ,.d_arid(split115_merge208_arid[(IDWID - 1):0])
    ,.d_arlen(split115_merge208_arlen[7:0])
    ,.d_arready(split115_merge208_arready)
    ,.d_arvalid(split115_merge208_arvalid)
    ,.d_awaddr(split115_merge208_awaddr[31:0])
    ,.d_awburst(split115_merge208_awburst[1:0])
    ,.d_awextras(split115_merge208_awextras[(EXTRAS - 1):0])
    ,.d_awid(split115_merge208_awid[(IDWID - 1):0])
    ,.d_awlen(split115_merge208_awlen[7:0])
    ,.d_awready(split115_merge208_awready)
    ,.d_awvalid(split115_merge208_awvalid)
    ,.d_bid(split115_merge208_bid[(IDWID - 1):0])
    ,.d_bready(split115_merge208_bready)
    ,.d_bresp(split115_merge208_bresp[1:0])
    ,.d_bvalid(split115_merge208_bvalid)
    ,.d_rdata(split115_merge208_rdata[(DWID - 1):0])
    ,.d_rid(split115_merge208_rid[(IDWID - 1):0])
    ,.d_rlast(split115_merge208_rlast)
    ,.d_rready(split115_merge208_rready)
    ,.d_rresp(split115_merge208_rresp[1:0])
    ,.d_rvalid(split115_merge208_rvalid)
    ,.d_wdata(split115_merge208_wdata[(DWID - 1):0])
    ,.d_wlast(split115_merge208_wlast)
    ,.d_wready(split115_merge208_wready)
    ,.d_wstrb(split115_merge208_wstrb[(WSTRB - 1):0])
    ,.d_wvalid(split115_merge208_wvalid)

);

axi_4_merger merge208 (
     .clk(clk),.rst_n(rst_n)
    ,.araddr(slv8_araddr[31:0])
    ,.arburst(slv8_arburst[1:0])
    ,.arextras(slv8_arextras[(EXTRAS - 1):0])
    ,.arid(slv8_arid[(IDWID - 1):0])
    ,.arlen(slv8_arlen[7:0])
    ,.arready(slv8_arready)
    ,.arvalid(slv8_arvalid)
    ,.awaddr(slv8_awaddr[31:0])
    ,.awburst(slv8_awburst[1:0])
    ,.awextras(slv8_awextras[(EXTRAS - 1):0])
    ,.awid(slv8_awid[3:0])
    ,.awlen(slv8_awlen[7:0])
    ,.awready(slv8_awready)
    ,.awvalid(slv8_awvalid)
    ,.bid(slv8_bid[(IDWID - 1):0])
    ,.bready(slv8_bready)
    ,.bresp(slv8_bresp[1:0])
    ,.bvalid(slv8_bvalid)
    ,.rid(slv8_rid[(IDWID - 1):0])
    ,.rlast(slv8_rlast)
    ,.rready(slv8_rready)
    ,.rresp(slv8_rresp[1:0])
    ,.rvalid(slv8_rvalid)
    ,.rdata(slv8_rdata[(DWID - 1):0])
    ,.wdata(slv8_wdata[(DWID - 1):0])
    ,.wlast(slv8_wlast)
    ,.wready(slv8_wready)
    ,.wstrb(slv8_wstrb[(WSTRB - 1):0])
    ,.wvalid(slv8_wvalid)


    ,.a_araddr(split100_merge208_araddr[31:0])
    ,.a_arburst(split100_merge208_arburst[1:0])
    ,.a_arextras(split100_merge208_arextras[(EXTRAS - 1):0])
    ,.a_arid(split100_merge208_arid[(IDWID - 1):0])
    ,.a_arlen(split100_merge208_arlen[7:0])
    ,.a_arready(split100_merge208_arready)
    ,.a_arvalid(split100_merge208_arvalid)
    ,.a_awaddr(split100_merge208_awaddr[31:0])
    ,.a_awburst(split100_merge208_awburst[1:0])
    ,.a_awextras(split100_merge208_awextras[(EXTRAS - 1):0])
    ,.a_awid(split100_merge208_awid[(IDWID - 1):0])
    ,.a_awlen(split100_merge208_awlen[7:0])
    ,.a_awready(split100_merge208_awready)
    ,.a_awvalid(split100_merge208_awvalid)
    ,.a_bid(split100_merge208_bid[(IDWID - 1):0])
    ,.a_bready(split100_merge208_bready)
    ,.a_bresp(split100_merge208_bresp[1:0])
    ,.a_bvalid(split100_merge208_bvalid)
    ,.a_rdata(split100_merge208_rdata[(DWID - 1):0])
    ,.a_rid(split100_merge208_rid[(IDWID - 1):0])
    ,.a_rlast(split100_merge208_rlast)
    ,.a_rready(split100_merge208_rready)
    ,.a_rresp(split100_merge208_rresp[1:0])
    ,.a_rvalid(split100_merge208_rvalid)
    ,.a_wdata(split100_merge208_wdata[(DWID - 1):0])
    ,.a_wlast(split100_merge208_wlast)
    ,.a_wready(split100_merge208_wready)
    ,.a_wstrb(split100_merge208_wstrb[(WSTRB - 1):0])
    ,.a_wvalid(split100_merge208_wvalid)

    ,.b_araddr(split105_merge208_araddr[31:0])
    ,.b_arburst(split105_merge208_arburst[1:0])
    ,.b_arextras(split105_merge208_arextras[(EXTRAS - 1):0])
    ,.b_arid(split105_merge208_arid[(IDWID - 1):0])
    ,.b_arlen(split105_merge208_arlen[7:0])
    ,.b_arready(split105_merge208_arready)
    ,.b_arvalid(split105_merge208_arvalid)
    ,.b_awaddr(split105_merge208_awaddr[31:0])
    ,.b_awburst(split105_merge208_awburst[1:0])
    ,.b_awextras(split105_merge208_awextras[(EXTRAS - 1):0])
    ,.b_awid(split105_merge208_awid[(IDWID - 1):0])
    ,.b_awlen(split105_merge208_awlen[7:0])
    ,.b_awready(split105_merge208_awready)
    ,.b_awvalid(split105_merge208_awvalid)
    ,.b_bid(split105_merge208_bid[(IDWID - 1):0])
    ,.b_bready(split105_merge208_bready)
    ,.b_bresp(split105_merge208_bresp[1:0])
    ,.b_bvalid(split105_merge208_bvalid)
    ,.b_rdata(split105_merge208_rdata[(DWID - 1):0])
    ,.b_rid(split105_merge208_rid[(IDWID - 1):0])
    ,.b_rlast(split105_merge208_rlast)
    ,.b_rready(split105_merge208_rready)
    ,.b_rresp(split105_merge208_rresp[1:0])
    ,.b_rvalid(split105_merge208_rvalid)
    ,.b_wdata(split105_merge208_wdata[(DWID - 1):0])
    ,.b_wlast(split105_merge208_wlast)
    ,.b_wready(split105_merge208_wready)
    ,.b_wstrb(split105_merge208_wstrb[(WSTRB - 1):0])
    ,.b_wvalid(split105_merge208_wvalid)

    ,.c_araddr(split114_merge208_araddr[31:0])
    ,.c_arburst(split114_merge208_arburst[1:0])
    ,.c_arextras(split114_merge208_arextras[(EXTRAS - 1):0])
    ,.c_arid(split114_merge208_arid[(IDWID - 1):0])
    ,.c_arlen(split114_merge208_arlen[7:0])
    ,.c_arready(split114_merge208_arready)
    ,.c_arvalid(split114_merge208_arvalid)
    ,.c_awaddr(split114_merge208_awaddr[31:0])
    ,.c_awburst(split114_merge208_awburst[1:0])
    ,.c_awextras(split114_merge208_awextras[(EXTRAS - 1):0])
    ,.c_awid(split114_merge208_awid[(IDWID - 1):0])
    ,.c_awlen(split114_merge208_awlen[7:0])
    ,.c_awready(split114_merge208_awready)
    ,.c_awvalid(split114_merge208_awvalid)
    ,.c_bid(split114_merge208_bid[(IDWID - 1):0])
    ,.c_bready(split114_merge208_bready)
    ,.c_bresp(split114_merge208_bresp[1:0])
    ,.c_bvalid(split114_merge208_bvalid)
    ,.c_rdata(split114_merge208_rdata[(DWID - 1):0])
    ,.c_rid(split114_merge208_rid[(IDWID - 1):0])
    ,.c_rlast(split114_merge208_rlast)
    ,.c_rready(split114_merge208_rready)
    ,.c_rresp(split114_merge208_rresp[1:0])
    ,.c_rvalid(split114_merge208_rvalid)
    ,.c_wdata(split114_merge208_wdata[(DWID - 1):0])
    ,.c_wlast(split114_merge208_wlast)
    ,.c_wready(split114_merge208_wready)
    ,.c_wstrb(split114_merge208_wstrb[(WSTRB - 1):0])
    ,.c_wvalid(split114_merge208_wvalid)

    ,.d_araddr(split115_merge208_araddr[31:0])
    ,.d_arburst(split115_merge208_arburst[1:0])
    ,.d_arextras(split115_merge208_arextras[(EXTRAS - 1):0])
    ,.d_arid(split115_merge208_arid[(IDWID - 1):0])
    ,.d_arlen(split115_merge208_arlen[7:0])
    ,.d_arready(split115_merge208_arready)
    ,.d_arvalid(split115_merge208_arvalid)
    ,.d_awaddr(split115_merge208_awaddr[31:0])
    ,.d_awburst(split115_merge208_awburst[1:0])
    ,.d_awextras(split115_merge208_awextras[(EXTRAS - 1):0])
    ,.d_awid(split115_merge208_awid[(IDWID - 1):0])
    ,.d_awlen(split115_merge208_awlen[7:0])
    ,.d_awready(split115_merge208_awready)
    ,.d_awvalid(split115_merge208_awvalid)
    ,.d_bid(split115_merge208_bid[(IDWID - 1):0])
    ,.d_bready(split115_merge208_bready)
    ,.d_bresp(split115_merge208_bresp[1:0])
    ,.d_bvalid(split115_merge208_bvalid)
    ,.d_rdata(split115_merge208_rdata[(DWID - 1):0])
    ,.d_rid(split115_merge208_rid[(IDWID - 1):0])
    ,.d_rlast(split115_merge208_rlast)
    ,.d_rready(split115_merge208_rready)
    ,.d_rresp(split115_merge208_rresp[1:0])
    ,.d_rvalid(split115_merge208_rvalid)
    ,.d_wdata(split115_merge208_wdata[(DWID - 1):0])
    ,.d_wlast(split115_merge208_wlast)
    ,.d_wready(split115_merge208_wready)
    ,.d_wstrb(split115_merge208_wstrb[(WSTRB - 1):0])
    ,.d_wvalid(split115_merge208_wvalid)
);


axi_4_merger merge211 (
     .clk(clk),.rst_n(rst_n)
    ,.araddr(slv11_araddr[31:0])
    ,.arburst(slv11_arburst[1:0])
    ,.arextras(slv11_arextras[(EXTRAS - 1):0])
    ,.arid(slv11_arid[(IDWID - 1):0])
    ,.arlen(slv11_arlen[7:0])
    ,.arready(slv11_arready)
    ,.arvalid(slv11_arvalid)
    ,.awaddr(slv11_awaddr[31:0])
    ,.awburst(slv11_awburst[1:0])
    ,.awextras(slv11_awextras[(EXTRAS - 1):0])
    ,.awid(slv11_awid[3:0])
    ,.awlen(slv11_awlen[7:0])
    ,.awready(slv11_awready)
    ,.awvalid(slv11_awvalid)
    ,.bid(slv11_bid[(IDWID - 1):0])
    ,.bready(slv11_bready)
    ,.bresp(slv11_bresp[1:0])
    ,.bvalid(slv11_bvalid)
    ,.rid(slv11_rid[(IDWID - 1):0])
    ,.rlast(slv11_rlast)
    ,.rready(slv11_rready)
    ,.rresp(slv11_rresp[1:0])
    ,.rvalid(slv11_rvalid)
    ,.rdata(slv11_rdata[(DWID - 1):0])
    ,.wdata(slv11_wdata[(DWID - 1):0])
    ,.wlast(slv11_wlast)
    ,.wready(slv11_wready)
    ,.wstrb(slv11_wstrb[(WSTRB - 1):0])
    ,.wvalid(slv11_wvalid)


    ,.a_araddr(split100_merge211_araddr[31:0])
    ,.a_arburst(split100_merge211_arburst[1:0])
    ,.a_arextras(split100_merge211_arextras[(EXTRAS - 1):0])
    ,.a_arid(split100_merge211_arid[(IDWID - 1):0])
    ,.a_arlen(split100_merge211_arlen[7:0])
    ,.a_arready(split100_merge211_arready)
    ,.a_arvalid(split100_merge211_arvalid)
    ,.a_awaddr(split100_merge211_awaddr[31:0])
    ,.a_awburst(split100_merge211_awburst[1:0])
    ,.a_awextras(split100_merge211_awextras[(EXTRAS - 1):0])
    ,.a_awid(split100_merge211_awid[(IDWID - 1):0])
    ,.a_awlen(split100_merge211_awlen[7:0])
    ,.a_awready(split100_merge211_awready)
    ,.a_awvalid(split100_merge211_awvalid)
    ,.a_bid(split100_merge211_bid[(IDWID - 1):0])
    ,.a_bready(split100_merge211_bready)
    ,.a_bresp(split100_merge211_bresp[1:0])
    ,.a_bvalid(split100_merge211_bvalid)
    ,.a_rdata(split100_merge211_rdata[(DWID - 1):0])
    ,.a_rid(split100_merge211_rid[(IDWID - 1):0])
    ,.a_rlast(split100_merge211_rlast)
    ,.a_rready(split100_merge211_rready)
    ,.a_rresp(split100_merge211_rresp[1:0])
    ,.a_rvalid(split100_merge211_rvalid)
    ,.a_wdata(split100_merge211_wdata[(DWID - 1):0])
    ,.a_wlast(split100_merge211_wlast)
    ,.a_wready(split100_merge211_wready)
    ,.a_wstrb(split100_merge211_wstrb[(WSTRB - 1):0])
    ,.a_wvalid(split100_merge211_wvalid)

    ,.b_araddr(split106_merge211_araddr[31:0])
    ,.b_arburst(split106_merge211_arburst[1:0])
    ,.b_arextras(split106_merge211_arextras[(EXTRAS - 1):0])
    ,.b_arid(split106_merge211_arid[(IDWID - 1):0])
    ,.b_arlen(split106_merge211_arlen[7:0])
    ,.b_arready(split106_merge211_arready)
    ,.b_arvalid(split106_merge211_arvalid)
    ,.b_awaddr(split106_merge211_awaddr[31:0])
    ,.b_awburst(split106_merge211_awburst[1:0])
    ,.b_awextras(split106_merge211_awextras[(EXTRAS - 1):0])
    ,.b_awid(split106_merge211_awid[(IDWID - 1):0])
    ,.b_awlen(split106_merge211_awlen[7:0])
    ,.b_awready(split106_merge211_awready)
    ,.b_awvalid(split106_merge211_awvalid)
    ,.b_bid(split106_merge211_bid[(IDWID - 1):0])
    ,.b_bready(split106_merge211_bready)
    ,.b_bresp(split106_merge211_bresp[1:0])
    ,.b_bvalid(split106_merge211_bvalid)
    ,.b_rdata(split106_merge211_rdata[(DWID - 1):0])
    ,.b_rid(split106_merge211_rid[(IDWID - 1):0])
    ,.b_rlast(split106_merge211_rlast)
    ,.b_rready(split106_merge211_rready)
    ,.b_rresp(split106_merge211_rresp[1:0])
    ,.b_rvalid(split106_merge211_rvalid)
    ,.b_wdata(split106_merge211_wdata[(DWID - 1):0])
    ,.b_wlast(split106_merge211_wlast)
    ,.b_wready(split106_merge211_wready)
    ,.b_wstrb(split106_merge211_wstrb[(WSTRB - 1):0])
    ,.b_wvalid(split106_merge211_wvalid)

    ,.c_araddr(split107_merge211_araddr[31:0])
    ,.c_arburst(split107_merge211_arburst[1:0])
    ,.c_arextras(split107_merge211_arextras[(EXTRAS - 1):0])
    ,.c_arid(split107_merge211_arid[(IDWID - 1):0])
    ,.c_arlen(split107_merge211_arlen[7:0])
    ,.c_arready(split107_merge211_arready)
    ,.c_arvalid(split107_merge211_arvalid)
    ,.c_awaddr(split107_merge211_awaddr[31:0])
    ,.c_awburst(split107_merge211_awburst[1:0])
    ,.c_awextras(split107_merge211_awextras[(EXTRAS - 1):0])
    ,.c_awid(split107_merge211_awid[(IDWID - 1):0])
    ,.c_awlen(split107_merge211_awlen[7:0])
    ,.c_awready(split107_merge211_awready)
    ,.c_awvalid(split107_merge211_awvalid)
    ,.c_bid(split107_merge211_bid[(IDWID - 1):0])
    ,.c_bready(split107_merge211_bready)
    ,.c_bresp(split107_merge211_bresp[1:0])
    ,.c_bvalid(split107_merge211_bvalid)
    ,.c_rdata(split107_merge211_rdata[(DWID - 1):0])
    ,.c_rid(split107_merge211_rid[(IDWID - 1):0])
    ,.c_rlast(split107_merge211_rlast)
    ,.c_rready(split107_merge211_rready)
    ,.c_rresp(split107_merge211_rresp[1:0])
    ,.c_rvalid(split107_merge211_rvalid)
    ,.c_wdata(split107_merge211_wdata[(DWID - 1):0])
    ,.c_wlast(split107_merge211_wlast)
    ,.c_wready(split107_merge211_wready)
    ,.c_wstrb(split107_merge211_wstrb[(WSTRB - 1):0])
    ,.c_wvalid(split107_merge211_wvalid)

    ,.d_araddr(split108_merge211_araddr[31:0])
    ,.d_arburst(split108_merge211_arburst[1:0])
    ,.d_arextras(split108_merge211_arextras[(EXTRAS - 1):0])
    ,.d_arid(split108_merge211_arid[(IDWID - 1):0])
    ,.d_arlen(split108_merge211_arlen[7:0])
    ,.d_arready(split108_merge211_arready)
    ,.d_arvalid(split108_merge211_arvalid)
    ,.d_awaddr(split108_merge211_awaddr[31:0])
    ,.d_awburst(split108_merge211_awburst[1:0])
    ,.d_awextras(split108_merge211_awextras[(EXTRAS - 1):0])
    ,.d_awid(split108_merge211_awid[(IDWID - 1):0])
    ,.d_awlen(split108_merge211_awlen[7:0])
    ,.d_awready(split108_merge211_awready)
    ,.d_awvalid(split108_merge211_awvalid)
    ,.d_bid(split108_merge211_bid[(IDWID - 1):0])
    ,.d_bready(split108_merge211_bready)
    ,.d_bresp(split108_merge211_bresp[1:0])
    ,.d_bvalid(split108_merge211_bvalid)
    ,.d_rdata(split108_merge211_rdata[(DWID - 1):0])
    ,.d_rid(split108_merge211_rid[(IDWID - 1):0])
    ,.d_rlast(split108_merge211_rlast)
    ,.d_rready(split108_merge211_rready)
    ,.d_rresp(split108_merge211_rresp[1:0])
    ,.d_rvalid(split108_merge211_rvalid)
    ,.d_wdata(split108_merge211_wdata[(DWID - 1):0])
    ,.d_wlast(split108_merge211_wlast)
    ,.d_wready(split108_merge211_wready)
    ,.d_wstrb(split108_merge211_wstrb[(WSTRB - 1):0])
    ,.d_wvalid(split108_merge211_wvalid)
);


axi_4_merger merge212 (
     .clk(clk),.rst_n(rst_n)
    ,.araddr(slv12_araddr[31:0])
    ,.arburst(slv12_arburst[1:0])
    ,.arextras(slv12_arextras[(EXTRAS - 1):0])
    ,.arid(slv12_arid[(IDWID - 1):0])
    ,.arlen(slv12_arlen[7:0])
    ,.arready(slv12_arready)
    ,.arvalid(slv12_arvalid)
    ,.awaddr(slv12_awaddr[31:0])
    ,.awburst(slv12_awburst[1:0])
    ,.awextras(slv12_awextras[(EXTRAS - 1):0])
    ,.awid(slv12_awid[3:0])
    ,.awlen(slv12_awlen[7:0])
    ,.awready(slv12_awready)
    ,.awvalid(slv12_awvalid)
    ,.bid(slv12_bid[(IDWID - 1):0])
    ,.bready(slv12_bready)
    ,.bresp(slv12_bresp[1:0])
    ,.bvalid(slv12_bvalid)
    ,.rid(slv12_rid[(IDWID - 1):0])
    ,.rlast(slv12_rlast)
    ,.rready(slv12_rready)
    ,.rresp(slv12_rresp[1:0])
    ,.rvalid(slv12_rvalid)
    ,.rdata(slv12_rdata[(DWID - 1):0])
    ,.wdata(slv12_wdata[(DWID - 1):0])
    ,.wlast(slv12_wlast)
    ,.wready(slv12_wready)
    ,.wstrb(slv12_wstrb[(WSTRB - 1):0])
    ,.wvalid(slv12_wvalid)


    ,.a_araddr(split100_merge212_araddr[31:0])
    ,.a_arburst(split100_merge212_arburst[1:0])
    ,.a_arextras(split100_merge212_arextras[(EXTRAS - 1):0])
    ,.a_arid(split100_merge212_arid[(IDWID - 1):0])
    ,.a_arlen(split100_merge212_arlen[7:0])
    ,.a_arready(split100_merge212_arready)
    ,.a_arvalid(split100_merge212_arvalid)
    ,.a_awaddr(split100_merge212_awaddr[31:0])
    ,.a_awburst(split100_merge212_awburst[1:0])
    ,.a_awextras(split100_merge212_awextras[(EXTRAS - 1):0])
    ,.a_awid(split100_merge212_awid[(IDWID - 1):0])
    ,.a_awlen(split100_merge212_awlen[7:0])
    ,.a_awready(split100_merge212_awready)
    ,.a_awvalid(split100_merge212_awvalid)
    ,.a_bid(split100_merge212_bid[(IDWID - 1):0])
    ,.a_bready(split100_merge212_bready)
    ,.a_bresp(split100_merge212_bresp[1:0])
    ,.a_bvalid(split100_merge212_bvalid)
    ,.a_rdata(split100_merge212_rdata[(DWID - 1):0])
    ,.a_rid(split100_merge212_rid[(IDWID - 1):0])
    ,.a_rlast(split100_merge212_rlast)
    ,.a_rready(split100_merge212_rready)
    ,.a_rresp(split100_merge212_rresp[1:0])
    ,.a_rvalid(split100_merge212_rvalid)
    ,.a_wdata(split100_merge212_wdata[(DWID - 1):0])
    ,.a_wlast(split100_merge212_wlast)
    ,.a_wready(split100_merge212_wready)
    ,.a_wstrb(split100_merge212_wstrb[(WSTRB - 1):0])
    ,.a_wvalid(split100_merge212_wvalid)

    ,.b_araddr(split101_merge212_araddr[31:0])
    ,.b_arburst(split101_merge212_arburst[1:0])
    ,.b_arextras(split101_merge212_arextras[(EXTRAS - 1):0])
    ,.b_arid(split101_merge212_arid[(IDWID - 1):0])
    ,.b_arlen(split101_merge212_arlen[7:0])
    ,.b_arready(split101_merge212_arready)
    ,.b_arvalid(split101_merge212_arvalid)
    ,.b_awaddr(split101_merge212_awaddr[31:0])
    ,.b_awburst(split101_merge212_awburst[1:0])
    ,.b_awextras(split101_merge212_awextras[(EXTRAS - 1):0])
    ,.b_awid(split101_merge212_awid[(IDWID - 1):0])
    ,.b_awlen(split101_merge212_awlen[7:0])
    ,.b_awready(split101_merge212_awready)
    ,.b_awvalid(split101_merge212_awvalid)
    ,.b_bid(split101_merge212_bid[(IDWID - 1):0])
    ,.b_bready(split101_merge212_bready)
    ,.b_bresp(split101_merge212_bresp[1:0])
    ,.b_bvalid(split101_merge212_bvalid)
    ,.b_rdata(split101_merge212_rdata[(DWID - 1):0])
    ,.b_rid(split101_merge212_rid[(IDWID - 1):0])
    ,.b_rlast(split101_merge212_rlast)
    ,.b_rready(split101_merge212_rready)
    ,.b_rresp(split101_merge212_rresp[1:0])
    ,.b_rvalid(split101_merge212_rvalid)
    ,.b_wdata(split101_merge212_wdata[(DWID - 1):0])
    ,.b_wlast(split101_merge212_wlast)
    ,.b_wready(split101_merge212_wready)
    ,.b_wstrb(split101_merge212_wstrb[(WSTRB - 1):0])
    ,.b_wvalid(split101_merge212_wvalid)

    ,.c_araddr(split105_merge212_araddr[31:0])
    ,.c_arburst(split105_merge212_arburst[1:0])
    ,.c_arextras(split105_merge212_arextras[(EXTRAS - 1):0])
    ,.c_arid(split105_merge212_arid[(IDWID - 1):0])
    ,.c_arlen(split105_merge212_arlen[7:0])
    ,.c_arready(split105_merge212_arready)
    ,.c_arvalid(split105_merge212_arvalid)
    ,.c_awaddr(split105_merge212_awaddr[31:0])
    ,.c_awburst(split105_merge212_awburst[1:0])
    ,.c_awextras(split105_merge212_awextras[(EXTRAS - 1):0])
    ,.c_awid(split105_merge212_awid[(IDWID - 1):0])
    ,.c_awlen(split105_merge212_awlen[7:0])
    ,.c_awready(split105_merge212_awready)
    ,.c_awvalid(split105_merge212_awvalid)
    ,.c_bid(split105_merge212_bid[(IDWID - 1):0])
    ,.c_bready(split105_merge212_bready)
    ,.c_bresp(split105_merge212_bresp[1:0])
    ,.c_bvalid(split105_merge212_bvalid)
    ,.c_rdata(split105_merge212_rdata[(DWID - 1):0])
    ,.c_rid(split105_merge212_rid[(IDWID - 1):0])
    ,.c_rlast(split105_merge212_rlast)
    ,.c_rready(split105_merge212_rready)
    ,.c_rresp(split105_merge212_rresp[1:0])
    ,.c_rvalid(split105_merge212_rvalid)
    ,.c_wdata(split105_merge212_wdata[(DWID - 1):0])
    ,.c_wlast(split105_merge212_wlast)
    ,.c_wready(split105_merge212_wready)
    ,.c_wstrb(split105_merge212_wstrb[(WSTRB - 1):0])
    ,.c_wvalid(split105_merge212_wvalid)

    ,.d_araddr(split113_merge212_araddr[31:0])
    ,.d_arburst(split113_merge212_arburst[1:0])
    ,.d_arextras(split113_merge212_arextras[(EXTRAS - 1):0])
    ,.d_arid(split113_merge212_arid[(IDWID - 1):0])
    ,.d_arlen(split113_merge212_arlen[7:0])
    ,.d_arready(split113_merge212_arready)
    ,.d_arvalid(split113_merge212_arvalid)
    ,.d_awaddr(split113_merge212_awaddr[31:0])
    ,.d_awburst(split113_merge212_awburst[1:0])
    ,.d_awextras(split113_merge212_awextras[(EXTRAS - 1):0])
    ,.d_awid(split113_merge212_awid[(IDWID - 1):0])
    ,.d_awlen(split113_merge212_awlen[7:0])
    ,.d_awready(split113_merge212_awready)
    ,.d_awvalid(split113_merge212_awvalid)
    ,.d_bid(split113_merge212_bid[(IDWID - 1):0])
    ,.d_bready(split113_merge212_bready)
    ,.d_bresp(split113_merge212_bresp[1:0])
    ,.d_bvalid(split113_merge212_bvalid)
    ,.d_rdata(split113_merge212_rdata[(DWID - 1):0])
    ,.d_rid(split113_merge212_rid[(IDWID - 1):0])
    ,.d_rlast(split113_merge212_rlast)
    ,.d_rready(split113_merge212_rready)
    ,.d_rresp(split113_merge212_rresp[1:0])
    ,.d_rvalid(split113_merge212_rvalid)
    ,.d_wdata(split113_merge212_wdata[(DWID - 1):0])
    ,.d_wlast(split113_merge212_wlast)
    ,.d_wready(split113_merge212_wready)
    ,.d_wstrb(split113_merge212_wstrb[(WSTRB - 1):0])
    ,.d_wvalid(split113_merge212_wvalid)
);


axi_4_merger merge206 (
     .clk(clk),.rst_n(rst_n)
    ,.araddr(slv6_araddr[31:0])
    ,.arburst(slv6_arburst[1:0])
    ,.arextras(slv6_arextras[(EXTRAS - 1):0])
    ,.arid(slv6_arid[(IDWID - 1):0])
    ,.arlen(slv6_arlen[7:0])
    ,.arready(slv6_arready)
    ,.arvalid(slv6_arvalid)
    ,.awaddr(slv6_awaddr[31:0])
    ,.awburst(slv6_awburst[1:0])
    ,.awextras(slv6_awextras[(EXTRAS - 1):0])
    ,.awid(slv6_awid[3:0])
    ,.awlen(slv6_awlen[7:0])
    ,.awready(slv6_awready)
    ,.awvalid(slv6_awvalid)
    ,.bid(slv6_bid[(IDWID - 1):0])
    ,.bready(slv6_bready)
    ,.bresp(slv6_bresp[1:0])
    ,.bvalid(slv6_bvalid)
    ,.rid(slv6_rid[(IDWID - 1):0])
    ,.rlast(slv6_rlast)
    ,.rready(slv6_rready)
    ,.rresp(slv6_rresp[1:0])
    ,.rvalid(slv6_rvalid)
    ,.rdata(slv6_rdata[(DWID - 1):0])
    ,.wdata(slv6_wdata[(DWID - 1):0])
    ,.wlast(slv6_wlast)
    ,.wready(slv6_wready)
    ,.wstrb(slv6_wstrb[(WSTRB - 1):0])
    ,.wvalid(slv6_wvalid)


    ,.a_araddr(split100_merge206_araddr[31:0])
    ,.a_arburst(split100_merge206_arburst[1:0])
    ,.a_arextras(split100_merge206_arextras[(EXTRAS - 1):0])
    ,.a_arid(split100_merge206_arid[(IDWID - 1):0])
    ,.a_arlen(split100_merge206_arlen[7:0])
    ,.a_arready(split100_merge206_arready)
    ,.a_arvalid(split100_merge206_arvalid)
    ,.a_awaddr(split100_merge206_awaddr[31:0])
    ,.a_awburst(split100_merge206_awburst[1:0])
    ,.a_awextras(split100_merge206_awextras[(EXTRAS - 1):0])
    ,.a_awid(split100_merge206_awid[(IDWID - 1):0])
    ,.a_awlen(split100_merge206_awlen[7:0])
    ,.a_awready(split100_merge206_awready)
    ,.a_awvalid(split100_merge206_awvalid)
    ,.a_bid(split100_merge206_bid[(IDWID - 1):0])
    ,.a_bready(split100_merge206_bready)
    ,.a_bresp(split100_merge206_bresp[1:0])
    ,.a_bvalid(split100_merge206_bvalid)
    ,.a_rdata(split100_merge206_rdata[(DWID - 1):0])
    ,.a_rid(split100_merge206_rid[(IDWID - 1):0])
    ,.a_rlast(split100_merge206_rlast)
    ,.a_rready(split100_merge206_rready)
    ,.a_rresp(split100_merge206_rresp[1:0])
    ,.a_rvalid(split100_merge206_rvalid)
    ,.a_wdata(split100_merge206_wdata[(DWID - 1):0])
    ,.a_wlast(split100_merge206_wlast)
    ,.a_wready(split100_merge206_wready)
    ,.a_wstrb(split100_merge206_wstrb[(WSTRB - 1):0])
    ,.a_wvalid(split100_merge206_wvalid)

    ,.b_araddr(split103_merge206_araddr[31:0])
    ,.b_arburst(split103_merge206_arburst[1:0])
    ,.b_arextras(split103_merge206_arextras[(EXTRAS - 1):0])
    ,.b_arid(split103_merge206_arid[(IDWID - 1):0])
    ,.b_arlen(split103_merge206_arlen[7:0])
    ,.b_arready(split103_merge206_arready)
    ,.b_arvalid(split103_merge206_arvalid)
    ,.b_awaddr(split103_merge206_awaddr[31:0])
    ,.b_awburst(split103_merge206_awburst[1:0])
    ,.b_awextras(split103_merge206_awextras[(EXTRAS - 1):0])
    ,.b_awid(split103_merge206_awid[(IDWID - 1):0])
    ,.b_awlen(split103_merge206_awlen[7:0])
    ,.b_awready(split103_merge206_awready)
    ,.b_awvalid(split103_merge206_awvalid)
    ,.b_bid(split103_merge206_bid[(IDWID - 1):0])
    ,.b_bready(split103_merge206_bready)
    ,.b_bresp(split103_merge206_bresp[1:0])
    ,.b_bvalid(split103_merge206_bvalid)
    ,.b_rdata(split103_merge206_rdata[(DWID - 1):0])
    ,.b_rid(split103_merge206_rid[(IDWID - 1):0])
    ,.b_rlast(split103_merge206_rlast)
    ,.b_rready(split103_merge206_rready)
    ,.b_rresp(split103_merge206_rresp[1:0])
    ,.b_rvalid(split103_merge206_rvalid)
    ,.b_wdata(split103_merge206_wdata[(DWID - 1):0])
    ,.b_wlast(split103_merge206_wlast)
    ,.b_wready(split103_merge206_wready)
    ,.b_wstrb(split103_merge206_wstrb[(WSTRB - 1):0])
    ,.b_wvalid(split103_merge206_wvalid)

    ,.c_araddr(split104_merge206_araddr[31:0])
    ,.c_arburst(split104_merge206_arburst[1:0])
    ,.c_arextras(split104_merge206_arextras[(EXTRAS - 1):0])
    ,.c_arid(split104_merge206_arid[(IDWID - 1):0])
    ,.c_arlen(split104_merge206_arlen[7:0])
    ,.c_arready(split104_merge206_arready)
    ,.c_arvalid(split104_merge206_arvalid)
    ,.c_awaddr(split104_merge206_awaddr[31:0])
    ,.c_awburst(split104_merge206_awburst[1:0])
    ,.c_awextras(split104_merge206_awextras[(EXTRAS - 1):0])
    ,.c_awid(split104_merge206_awid[(IDWID - 1):0])
    ,.c_awlen(split104_merge206_awlen[7:0])
    ,.c_awready(split104_merge206_awready)
    ,.c_awvalid(split104_merge206_awvalid)
    ,.c_bid(split104_merge206_bid[(IDWID - 1):0])
    ,.c_bready(split104_merge206_bready)
    ,.c_bresp(split104_merge206_bresp[1:0])
    ,.c_bvalid(split104_merge206_bvalid)
    ,.c_rdata(split104_merge206_rdata[(DWID - 1):0])
    ,.c_rid(split104_merge206_rid[(IDWID - 1):0])
    ,.c_rlast(split104_merge206_rlast)
    ,.c_rready(split104_merge206_rready)
    ,.c_rresp(split104_merge206_rresp[1:0])
    ,.c_rvalid(split104_merge206_rvalid)
    ,.c_wdata(split104_merge206_wdata[(DWID - 1):0])
    ,.c_wlast(split104_merge206_wlast)
    ,.c_wready(split104_merge206_wready)
    ,.c_wstrb(split104_merge206_wstrb[(WSTRB - 1):0])
    ,.c_wvalid(split104_merge206_wvalid)

    ,.d_araddr(split113_merge206_araddr[31:0])
    ,.d_arburst(split113_merge206_arburst[1:0])
    ,.d_arextras(split113_merge206_arextras[(EXTRAS - 1):0])
    ,.d_arid(split113_merge206_arid[(IDWID - 1):0])
    ,.d_arlen(split113_merge206_arlen[7:0])
    ,.d_arready(split113_merge206_arready)
    ,.d_arvalid(split113_merge206_arvalid)
    ,.d_awaddr(split113_merge206_awaddr[31:0])
    ,.d_awburst(split113_merge206_awburst[1:0])
    ,.d_awextras(split113_merge206_awextras[(EXTRAS - 1):0])
    ,.d_awid(split113_merge206_awid[(IDWID - 1):0])
    ,.d_awlen(split113_merge206_awlen[7:0])
    ,.d_awready(split113_merge206_awready)
    ,.d_awvalid(split113_merge206_awvalid)
    ,.d_bid(split113_merge206_bid[(IDWID - 1):0])
    ,.d_bready(split113_merge206_bready)
    ,.d_bresp(split113_merge206_bresp[1:0])
    ,.d_bvalid(split113_merge206_bvalid)
    ,.d_rdata(split113_merge206_rdata[(DWID - 1):0])
    ,.d_rid(split113_merge206_rid[(IDWID - 1):0])
    ,.d_rlast(split113_merge206_rlast)
    ,.d_rready(split113_merge206_rready)
    ,.d_rresp(split113_merge206_rresp[1:0])
    ,.d_rvalid(split113_merge206_rvalid)
    ,.d_wdata(split113_merge206_wdata[(DWID - 1):0])
    ,.d_wlast(split113_merge206_wlast)
    ,.d_wready(split113_merge206_wready)
    ,.d_wstrb(split113_merge206_wstrb[(WSTRB - 1):0])
    ,.d_wvalid(split113_merge206_wvalid)
);


axi_4_merger merge203 (
     .clk(clk),.rst_n(rst_n)
    ,.araddr(slv3_araddr[31:0])
    ,.arburst(slv3_arburst[1:0])
    ,.arextras(slv3_arextras[(EXTRAS - 1):0])
    ,.arid(slv3_arid[(IDWID - 1):0])
    ,.arlen(slv3_arlen[7:0])
    ,.arready(slv3_arready)
    ,.arvalid(slv3_arvalid)
    ,.awaddr(slv3_awaddr[31:0])
    ,.awburst(slv3_awburst[1:0])
    ,.awextras(slv3_awextras[(EXTRAS - 1):0])
    ,.awid(slv3_awid[3:0])
    ,.awlen(slv3_awlen[7:0])
    ,.awready(slv3_awready)
    ,.awvalid(slv3_awvalid)
    ,.bid(slv3_bid[(IDWID - 1):0])
    ,.bready(slv3_bready)
    ,.bresp(slv3_bresp[1:0])
    ,.bvalid(slv3_bvalid)
    ,.rid(slv3_rid[(IDWID - 1):0])
    ,.rlast(slv3_rlast)
    ,.rready(slv3_rready)
    ,.rresp(slv3_rresp[1:0])
    ,.rvalid(slv3_rvalid)
    ,.rdata(slv3_rdata[(DWID - 1):0])
    ,.wdata(slv3_wdata[(DWID - 1):0])
    ,.wlast(slv3_wlast)
    ,.wready(slv3_wready)
    ,.wstrb(slv3_wstrb[(WSTRB - 1):0])
    ,.wvalid(slv3_wvalid)


    ,.a_araddr(split101_merge203_araddr[31:0])
    ,.a_arburst(split101_merge203_arburst[1:0])
    ,.a_arextras(split101_merge203_arextras[(EXTRAS - 1):0])
    ,.a_arid(split101_merge203_arid[(IDWID - 1):0])
    ,.a_arlen(split101_merge203_arlen[7:0])
    ,.a_arready(split101_merge203_arready)
    ,.a_arvalid(split101_merge203_arvalid)
    ,.a_awaddr(split101_merge203_awaddr[31:0])
    ,.a_awburst(split101_merge203_awburst[1:0])
    ,.a_awextras(split101_merge203_awextras[(EXTRAS - 1):0])
    ,.a_awid(split101_merge203_awid[(IDWID - 1):0])
    ,.a_awlen(split101_merge203_awlen[7:0])
    ,.a_awready(split101_merge203_awready)
    ,.a_awvalid(split101_merge203_awvalid)
    ,.a_bid(split101_merge203_bid[(IDWID - 1):0])
    ,.a_bready(split101_merge203_bready)
    ,.a_bresp(split101_merge203_bresp[1:0])
    ,.a_bvalid(split101_merge203_bvalid)
    ,.a_rdata(split101_merge203_rdata[(DWID - 1):0])
    ,.a_rid(split101_merge203_rid[(IDWID - 1):0])
    ,.a_rlast(split101_merge203_rlast)
    ,.a_rready(split101_merge203_rready)
    ,.a_rresp(split101_merge203_rresp[1:0])
    ,.a_rvalid(split101_merge203_rvalid)
    ,.a_wdata(split101_merge203_wdata[(DWID - 1):0])
    ,.a_wlast(split101_merge203_wlast)
    ,.a_wready(split101_merge203_wready)
    ,.a_wstrb(split101_merge203_wstrb[(WSTRB - 1):0])
    ,.a_wvalid(split101_merge203_wvalid)

    ,.b_araddr(split103_merge203_araddr[31:0])
    ,.b_arburst(split103_merge203_arburst[1:0])
    ,.b_arextras(split103_merge203_arextras[(EXTRAS - 1):0])
    ,.b_arid(split103_merge203_arid[(IDWID - 1):0])
    ,.b_arlen(split103_merge203_arlen[7:0])
    ,.b_arready(split103_merge203_arready)
    ,.b_arvalid(split103_merge203_arvalid)
    ,.b_awaddr(split103_merge203_awaddr[31:0])
    ,.b_awburst(split103_merge203_awburst[1:0])
    ,.b_awextras(split103_merge203_awextras[(EXTRAS - 1):0])
    ,.b_awid(split103_merge203_awid[(IDWID - 1):0])
    ,.b_awlen(split103_merge203_awlen[7:0])
    ,.b_awready(split103_merge203_awready)
    ,.b_awvalid(split103_merge203_awvalid)
    ,.b_bid(split103_merge203_bid[(IDWID - 1):0])
    ,.b_bready(split103_merge203_bready)
    ,.b_bresp(split103_merge203_bresp[1:0])
    ,.b_bvalid(split103_merge203_bvalid)
    ,.b_rdata(split103_merge203_rdata[(DWID - 1):0])
    ,.b_rid(split103_merge203_rid[(IDWID - 1):0])
    ,.b_rlast(split103_merge203_rlast)
    ,.b_rready(split103_merge203_rready)
    ,.b_rresp(split103_merge203_rresp[1:0])
    ,.b_rvalid(split103_merge203_rvalid)
    ,.b_wdata(split103_merge203_wdata[(DWID - 1):0])
    ,.b_wlast(split103_merge203_wlast)
    ,.b_wready(split103_merge203_wready)
    ,.b_wstrb(split103_merge203_wstrb[(WSTRB - 1):0])
    ,.b_wvalid(split103_merge203_wvalid)

    ,.c_araddr(split109_merge203_araddr[31:0])
    ,.c_arburst(split109_merge203_arburst[1:0])
    ,.c_arextras(split109_merge203_arextras[(EXTRAS - 1):0])
    ,.c_arid(split109_merge203_arid[(IDWID - 1):0])
    ,.c_arlen(split109_merge203_arlen[7:0])
    ,.c_arready(split109_merge203_arready)
    ,.c_arvalid(split109_merge203_arvalid)
    ,.c_awaddr(split109_merge203_awaddr[31:0])
    ,.c_awburst(split109_merge203_awburst[1:0])
    ,.c_awextras(split109_merge203_awextras[(EXTRAS - 1):0])
    ,.c_awid(split109_merge203_awid[(IDWID - 1):0])
    ,.c_awlen(split109_merge203_awlen[7:0])
    ,.c_awready(split109_merge203_awready)
    ,.c_awvalid(split109_merge203_awvalid)
    ,.c_bid(split109_merge203_bid[(IDWID - 1):0])
    ,.c_bready(split109_merge203_bready)
    ,.c_bresp(split109_merge203_bresp[1:0])
    ,.c_bvalid(split109_merge203_bvalid)
    ,.c_rdata(split109_merge203_rdata[(DWID - 1):0])
    ,.c_rid(split109_merge203_rid[(IDWID - 1):0])
    ,.c_rlast(split109_merge203_rlast)
    ,.c_rready(split109_merge203_rready)
    ,.c_rresp(split109_merge203_rresp[1:0])
    ,.c_rvalid(split109_merge203_rvalid)
    ,.c_wdata(split109_merge203_wdata[(DWID - 1):0])
    ,.c_wlast(split109_merge203_wlast)
    ,.c_wready(split109_merge203_wready)
    ,.c_wstrb(split109_merge203_wstrb[(WSTRB - 1):0])
    ,.c_wvalid(split109_merge203_wvalid)

    ,.d_araddr(split110_merge203_araddr[31:0])
    ,.d_arburst(split110_merge203_arburst[1:0])
    ,.d_arextras(split110_merge203_arextras[(EXTRAS - 1):0])
    ,.d_arid(split110_merge203_arid[(IDWID - 1):0])
    ,.d_arlen(split110_merge203_arlen[7:0])
    ,.d_arready(split110_merge203_arready)
    ,.d_arvalid(split110_merge203_arvalid)
    ,.d_awaddr(split110_merge203_awaddr[31:0])
    ,.d_awburst(split110_merge203_awburst[1:0])
    ,.d_awextras(split110_merge203_awextras[(EXTRAS - 1):0])
    ,.d_awid(split110_merge203_awid[(IDWID - 1):0])
    ,.d_awlen(split110_merge203_awlen[7:0])
    ,.d_awready(split110_merge203_awready)
    ,.d_awvalid(split110_merge203_awvalid)
    ,.d_bid(split110_merge203_bid[(IDWID - 1):0])
    ,.d_bready(split110_merge203_bready)
    ,.d_bresp(split110_merge203_bresp[1:0])
    ,.d_bvalid(split110_merge203_bvalid)
    ,.d_rdata(split110_merge203_rdata[(DWID - 1):0])
    ,.d_rid(split110_merge203_rid[(IDWID - 1):0])
    ,.d_rlast(split110_merge203_rlast)
    ,.d_rready(split110_merge203_rready)
    ,.d_rresp(split110_merge203_rresp[1:0])
    ,.d_rvalid(split110_merge203_rvalid)
    ,.d_wdata(split110_merge203_wdata[(DWID - 1):0])
    ,.d_wlast(split110_merge203_wlast)
    ,.d_wready(split110_merge203_wready)
    ,.d_wstrb(split110_merge203_wstrb[(WSTRB - 1):0])
    ,.d_wvalid(split110_merge203_wvalid)
);


axi_4_merger merge201 (
     .clk(clk),.rst_n(rst_n)
    ,.araddr(slv1_araddr[31:0])
    ,.arburst(slv1_arburst[1:0])
    ,.arextras(slv1_arextras[(EXTRAS - 1):0])
    ,.arid(slv1_arid[(IDWID - 1):0])
    ,.arlen(slv1_arlen[7:0])
    ,.arready(slv1_arready)
    ,.arvalid(slv1_arvalid)
    ,.awaddr(slv1_awaddr[31:0])
    ,.awburst(slv1_awburst[1:0])
    ,.awextras(slv1_awextras[(EXTRAS - 1):0])
    ,.awid(slv1_awid[3:0])
    ,.awlen(slv1_awlen[7:0])
    ,.awready(slv1_awready)
    ,.awvalid(slv1_awvalid)
    ,.bid(slv1_bid[(IDWID - 1):0])
    ,.bready(slv1_bready)
    ,.bresp(slv1_bresp[1:0])
    ,.bvalid(slv1_bvalid)
    ,.rid(slv1_rid[(IDWID - 1):0])
    ,.rlast(slv1_rlast)
    ,.rready(slv1_rready)
    ,.rresp(slv1_rresp[1:0])
    ,.rvalid(slv1_rvalid)
    ,.rdata(slv1_rdata[(DWID - 1):0])
    ,.wdata(slv1_wdata[(DWID - 1):0])
    ,.wlast(slv1_wlast)
    ,.wready(slv1_wready)
    ,.wstrb(slv1_wstrb[(WSTRB - 1):0])
    ,.wvalid(slv1_wvalid)


    ,.a_araddr(split101_merge201_araddr[31:0])
    ,.a_arburst(split101_merge201_arburst[1:0])
    ,.a_arextras(split101_merge201_arextras[(EXTRAS - 1):0])
    ,.a_arid(split101_merge201_arid[(IDWID - 1):0])
    ,.a_arlen(split101_merge201_arlen[7:0])
    ,.a_arready(split101_merge201_arready)
    ,.a_arvalid(split101_merge201_arvalid)
    ,.a_awaddr(split101_merge201_awaddr[31:0])
    ,.a_awburst(split101_merge201_awburst[1:0])
    ,.a_awextras(split101_merge201_awextras[(EXTRAS - 1):0])
    ,.a_awid(split101_merge201_awid[(IDWID - 1):0])
    ,.a_awlen(split101_merge201_awlen[7:0])
    ,.a_awready(split101_merge201_awready)
    ,.a_awvalid(split101_merge201_awvalid)
    ,.a_bid(split101_merge201_bid[(IDWID - 1):0])
    ,.a_bready(split101_merge201_bready)
    ,.a_bresp(split101_merge201_bresp[1:0])
    ,.a_bvalid(split101_merge201_bvalid)
    ,.a_rdata(split101_merge201_rdata[(DWID - 1):0])
    ,.a_rid(split101_merge201_rid[(IDWID - 1):0])
    ,.a_rlast(split101_merge201_rlast)
    ,.a_rready(split101_merge201_rready)
    ,.a_rresp(split101_merge201_rresp[1:0])
    ,.a_rvalid(split101_merge201_rvalid)
    ,.a_wdata(split101_merge201_wdata[(DWID - 1):0])
    ,.a_wlast(split101_merge201_wlast)
    ,.a_wready(split101_merge201_wready)
    ,.a_wstrb(split101_merge201_wstrb[(WSTRB - 1):0])
    ,.a_wvalid(split101_merge201_wvalid)

    ,.b_araddr(split102_merge201_araddr[31:0])
    ,.b_arburst(split102_merge201_arburst[1:0])
    ,.b_arextras(split102_merge201_arextras[(EXTRAS - 1):0])
    ,.b_arid(split102_merge201_arid[(IDWID - 1):0])
    ,.b_arlen(split102_merge201_arlen[7:0])
    ,.b_arready(split102_merge201_arready)
    ,.b_arvalid(split102_merge201_arvalid)
    ,.b_awaddr(split102_merge201_awaddr[31:0])
    ,.b_awburst(split102_merge201_awburst[1:0])
    ,.b_awextras(split102_merge201_awextras[(EXTRAS - 1):0])
    ,.b_awid(split102_merge201_awid[(IDWID - 1):0])
    ,.b_awlen(split102_merge201_awlen[7:0])
    ,.b_awready(split102_merge201_awready)
    ,.b_awvalid(split102_merge201_awvalid)
    ,.b_bid(split102_merge201_bid[(IDWID - 1):0])
    ,.b_bready(split102_merge201_bready)
    ,.b_bresp(split102_merge201_bresp[1:0])
    ,.b_bvalid(split102_merge201_bvalid)
    ,.b_rdata(split102_merge201_rdata[(DWID - 1):0])
    ,.b_rid(split102_merge201_rid[(IDWID - 1):0])
    ,.b_rlast(split102_merge201_rlast)
    ,.b_rready(split102_merge201_rready)
    ,.b_rresp(split102_merge201_rresp[1:0])
    ,.b_rvalid(split102_merge201_rvalid)
    ,.b_wdata(split102_merge201_wdata[(DWID - 1):0])
    ,.b_wlast(split102_merge201_wlast)
    ,.b_wready(split102_merge201_wready)
    ,.b_wstrb(split102_merge201_wstrb[(WSTRB - 1):0])
    ,.b_wvalid(split102_merge201_wvalid)

    ,.c_araddr(split112_merge201_araddr[31:0])
    ,.c_arburst(split112_merge201_arburst[1:0])
    ,.c_arextras(split112_merge201_arextras[(EXTRAS - 1):0])
    ,.c_arid(split112_merge201_arid[(IDWID - 1):0])
    ,.c_arlen(split112_merge201_arlen[7:0])
    ,.c_arready(split112_merge201_arready)
    ,.c_arvalid(split112_merge201_arvalid)
    ,.c_awaddr(split112_merge201_awaddr[31:0])
    ,.c_awburst(split112_merge201_awburst[1:0])
    ,.c_awextras(split112_merge201_awextras[(EXTRAS - 1):0])
    ,.c_awid(split112_merge201_awid[(IDWID - 1):0])
    ,.c_awlen(split112_merge201_awlen[7:0])
    ,.c_awready(split112_merge201_awready)
    ,.c_awvalid(split112_merge201_awvalid)
    ,.c_bid(split112_merge201_bid[(IDWID - 1):0])
    ,.c_bready(split112_merge201_bready)
    ,.c_bresp(split112_merge201_bresp[1:0])
    ,.c_bvalid(split112_merge201_bvalid)
    ,.c_rdata(split112_merge201_rdata[(DWID - 1):0])
    ,.c_rid(split112_merge201_rid[(IDWID - 1):0])
    ,.c_rlast(split112_merge201_rlast)
    ,.c_rready(split112_merge201_rready)
    ,.c_rresp(split112_merge201_rresp[1:0])
    ,.c_rvalid(split112_merge201_rvalid)
    ,.c_wdata(split112_merge201_wdata[(DWID - 1):0])
    ,.c_wlast(split112_merge201_wlast)
    ,.c_wready(split112_merge201_wready)
    ,.c_wstrb(split112_merge201_wstrb[(WSTRB - 1):0])
    ,.c_wvalid(split112_merge201_wvalid)

    ,.d_araddr(split113_merge201_araddr[31:0])
    ,.d_arburst(split113_merge201_arburst[1:0])
    ,.d_arextras(split113_merge201_arextras[(EXTRAS - 1):0])
    ,.d_arid(split113_merge201_arid[(IDWID - 1):0])
    ,.d_arlen(split113_merge201_arlen[7:0])
    ,.d_arready(split113_merge201_arready)
    ,.d_arvalid(split113_merge201_arvalid)
    ,.d_awaddr(split113_merge201_awaddr[31:0])
    ,.d_awburst(split113_merge201_awburst[1:0])
    ,.d_awextras(split113_merge201_awextras[(EXTRAS - 1):0])
    ,.d_awid(split113_merge201_awid[(IDWID - 1):0])
    ,.d_awlen(split113_merge201_awlen[7:0])
    ,.d_awready(split113_merge201_awready)
    ,.d_awvalid(split113_merge201_awvalid)
    ,.d_bid(split113_merge201_bid[(IDWID - 1):0])
    ,.d_bready(split113_merge201_bready)
    ,.d_bresp(split113_merge201_bresp[1:0])
    ,.d_bvalid(split113_merge201_bvalid)
    ,.d_rdata(split113_merge201_rdata[(DWID - 1):0])
    ,.d_rid(split113_merge201_rid[(IDWID - 1):0])
    ,.d_rlast(split113_merge201_rlast)
    ,.d_rready(split113_merge201_rready)
    ,.d_rresp(split113_merge201_rresp[1:0])
    ,.d_rvalid(split113_merge201_rvalid)
    ,.d_wdata(split113_merge201_wdata[(DWID - 1):0])
    ,.d_wlast(split113_merge201_wlast)
    ,.d_wready(split113_merge201_wready)
    ,.d_wstrb(split113_merge201_wstrb[(WSTRB - 1):0])
    ,.d_wvalid(split113_merge201_wvalid)
);


axi_4_merger merge209 (
     .clk(clk),.rst_n(rst_n)
    ,.araddr(slv9_araddr[31:0])
    ,.arburst(slv9_arburst[1:0])
    ,.arextras(slv9_arextras[(EXTRAS - 1):0])
    ,.arid(slv9_arid[(IDWID - 1):0])
    ,.arlen(slv9_arlen[7:0])
    ,.arready(slv9_arready)
    ,.arvalid(slv9_arvalid)
    ,.awaddr(slv9_awaddr[31:0])
    ,.awburst(slv9_awburst[1:0])
    ,.awextras(slv9_awextras[(EXTRAS - 1):0])
    ,.awid(slv9_awid[3:0])
    ,.awlen(slv9_awlen[7:0])
    ,.awready(slv9_awready)
    ,.awvalid(slv9_awvalid)
    ,.bid(slv9_bid[(IDWID - 1):0])
    ,.bready(slv9_bready)
    ,.bresp(slv9_bresp[1:0])
    ,.bvalid(slv9_bvalid)
    ,.rid(slv9_rid[(IDWID - 1):0])
    ,.rlast(slv9_rlast)
    ,.rready(slv9_rready)
    ,.rresp(slv9_rresp[1:0])
    ,.rvalid(slv9_rvalid)
    ,.rdata(slv9_rdata[(DWID - 1):0])
    ,.wdata(slv9_wdata[(DWID - 1):0])
    ,.wlast(slv9_wlast)
    ,.wready(slv9_wready)
    ,.wstrb(slv9_wstrb[(WSTRB - 1):0])
    ,.wvalid(slv9_wvalid)


    ,.a_araddr(split101_merge209_araddr[31:0])
    ,.a_arburst(split101_merge209_arburst[1:0])
    ,.a_arextras(split101_merge209_arextras[(EXTRAS - 1):0])
    ,.a_arid(split101_merge209_arid[(IDWID - 1):0])
    ,.a_arlen(split101_merge209_arlen[7:0])
    ,.a_arready(split101_merge209_arready)
    ,.a_arvalid(split101_merge209_arvalid)
    ,.a_awaddr(split101_merge209_awaddr[31:0])
    ,.a_awburst(split101_merge209_awburst[1:0])
    ,.a_awextras(split101_merge209_awextras[(EXTRAS - 1):0])
    ,.a_awid(split101_merge209_awid[(IDWID - 1):0])
    ,.a_awlen(split101_merge209_awlen[7:0])
    ,.a_awready(split101_merge209_awready)
    ,.a_awvalid(split101_merge209_awvalid)
    ,.a_bid(split101_merge209_bid[(IDWID - 1):0])
    ,.a_bready(split101_merge209_bready)
    ,.a_bresp(split101_merge209_bresp[1:0])
    ,.a_bvalid(split101_merge209_bvalid)
    ,.a_rdata(split101_merge209_rdata[(DWID - 1):0])
    ,.a_rid(split101_merge209_rid[(IDWID - 1):0])
    ,.a_rlast(split101_merge209_rlast)
    ,.a_rready(split101_merge209_rready)
    ,.a_rresp(split101_merge209_rresp[1:0])
    ,.a_rvalid(split101_merge209_rvalid)
    ,.a_wdata(split101_merge209_wdata[(DWID - 1):0])
    ,.a_wlast(split101_merge209_wlast)
    ,.a_wready(split101_merge209_wready)
    ,.a_wstrb(split101_merge209_wstrb[(WSTRB - 1):0])
    ,.a_wvalid(split101_merge209_wvalid)

    ,.b_araddr(split104_merge209_araddr[31:0])
    ,.b_arburst(split104_merge209_arburst[1:0])
    ,.b_arextras(split104_merge209_arextras[(EXTRAS - 1):0])
    ,.b_arid(split104_merge209_arid[(IDWID - 1):0])
    ,.b_arlen(split104_merge209_arlen[7:0])
    ,.b_arready(split104_merge209_arready)
    ,.b_arvalid(split104_merge209_arvalid)
    ,.b_awaddr(split104_merge209_awaddr[31:0])
    ,.b_awburst(split104_merge209_awburst[1:0])
    ,.b_awextras(split104_merge209_awextras[(EXTRAS - 1):0])
    ,.b_awid(split104_merge209_awid[(IDWID - 1):0])
    ,.b_awlen(split104_merge209_awlen[7:0])
    ,.b_awready(split104_merge209_awready)
    ,.b_awvalid(split104_merge209_awvalid)
    ,.b_bid(split104_merge209_bid[(IDWID - 1):0])
    ,.b_bready(split104_merge209_bready)
    ,.b_bresp(split104_merge209_bresp[1:0])
    ,.b_bvalid(split104_merge209_bvalid)
    ,.b_rdata(split104_merge209_rdata[(DWID - 1):0])
    ,.b_rid(split104_merge209_rid[(IDWID - 1):0])
    ,.b_rlast(split104_merge209_rlast)
    ,.b_rready(split104_merge209_rready)
    ,.b_rresp(split104_merge209_rresp[1:0])
    ,.b_rvalid(split104_merge209_rvalid)
    ,.b_wdata(split104_merge209_wdata[(DWID - 1):0])
    ,.b_wlast(split104_merge209_wlast)
    ,.b_wready(split104_merge209_wready)
    ,.b_wstrb(split104_merge209_wstrb[(WSTRB - 1):0])
    ,.b_wvalid(split104_merge209_wvalid)

    ,.c_araddr(split109_merge209_araddr[31:0])
    ,.c_arburst(split109_merge209_arburst[1:0])
    ,.c_arextras(split109_merge209_arextras[(EXTRAS - 1):0])
    ,.c_arid(split109_merge209_arid[(IDWID - 1):0])
    ,.c_arlen(split109_merge209_arlen[7:0])
    ,.c_arready(split109_merge209_arready)
    ,.c_arvalid(split109_merge209_arvalid)
    ,.c_awaddr(split109_merge209_awaddr[31:0])
    ,.c_awburst(split109_merge209_awburst[1:0])
    ,.c_awextras(split109_merge209_awextras[(EXTRAS - 1):0])
    ,.c_awid(split109_merge209_awid[(IDWID - 1):0])
    ,.c_awlen(split109_merge209_awlen[7:0])
    ,.c_awready(split109_merge209_awready)
    ,.c_awvalid(split109_merge209_awvalid)
    ,.c_bid(split109_merge209_bid[(IDWID - 1):0])
    ,.c_bready(split109_merge209_bready)
    ,.c_bresp(split109_merge209_bresp[1:0])
    ,.c_bvalid(split109_merge209_bvalid)
    ,.c_rdata(split109_merge209_rdata[(DWID - 1):0])
    ,.c_rid(split109_merge209_rid[(IDWID - 1):0])
    ,.c_rlast(split109_merge209_rlast)
    ,.c_rready(split109_merge209_rready)
    ,.c_rresp(split109_merge209_rresp[1:0])
    ,.c_rvalid(split109_merge209_rvalid)
    ,.c_wdata(split109_merge209_wdata[(DWID - 1):0])
    ,.c_wlast(split109_merge209_wlast)
    ,.c_wready(split109_merge209_wready)
    ,.c_wstrb(split109_merge209_wstrb[(WSTRB - 1):0])
    ,.c_wvalid(split109_merge209_wvalid)

    ,.d_araddr(split110_merge209_araddr[31:0])
    ,.d_arburst(split110_merge209_arburst[1:0])
    ,.d_arextras(split110_merge209_arextras[(EXTRAS - 1):0])
    ,.d_arid(split110_merge209_arid[(IDWID - 1):0])
    ,.d_arlen(split110_merge209_arlen[7:0])
    ,.d_arready(split110_merge209_arready)
    ,.d_arvalid(split110_merge209_arvalid)
    ,.d_awaddr(split110_merge209_awaddr[31:0])
    ,.d_awburst(split110_merge209_awburst[1:0])
    ,.d_awextras(split110_merge209_awextras[(EXTRAS - 1):0])
    ,.d_awid(split110_merge209_awid[(IDWID - 1):0])
    ,.d_awlen(split110_merge209_awlen[7:0])
    ,.d_awready(split110_merge209_awready)
    ,.d_awvalid(split110_merge209_awvalid)
    ,.d_bid(split110_merge209_bid[(IDWID - 1):0])
    ,.d_bready(split110_merge209_bready)
    ,.d_bresp(split110_merge209_bresp[1:0])
    ,.d_bvalid(split110_merge209_bvalid)
    ,.d_rdata(split110_merge209_rdata[(DWID - 1):0])
    ,.d_rid(split110_merge209_rid[(IDWID - 1):0])
    ,.d_rlast(split110_merge209_rlast)
    ,.d_rready(split110_merge209_rready)
    ,.d_rresp(split110_merge209_rresp[1:0])
    ,.d_rvalid(split110_merge209_rvalid)
    ,.d_wdata(split110_merge209_wdata[(DWID - 1):0])
    ,.d_wlast(split110_merge209_wlast)
    ,.d_wready(split110_merge209_wready)
    ,.d_wstrb(split110_merge209_wstrb[(WSTRB - 1):0])
    ,.d_wvalid(split110_merge209_wvalid)
);


axi_4_merger merge200 (
     .clk(clk),.rst_n(rst_n)
    ,.araddr(slv0_araddr[31:0])
    ,.arburst(slv0_arburst[1:0])
    ,.arextras(slv0_arextras[(EXTRAS - 1):0])
    ,.arid(slv0_arid[(IDWID - 1):0])
    ,.arlen(slv0_arlen[7:0])
    ,.arready(slv0_arready)
    ,.arvalid(slv0_arvalid)
    ,.awaddr(slv0_awaddr[31:0])
    ,.awburst(slv0_awburst[1:0])
    ,.awextras(slv0_awextras[(EXTRAS - 1):0])
    ,.awid(slv0_awid[3:0])
    ,.awlen(slv0_awlen[7:0])
    ,.awready(slv0_awready)
    ,.awvalid(slv0_awvalid)
    ,.bid(slv0_bid[(IDWID - 1):0])
    ,.bready(slv0_bready)
    ,.bresp(slv0_bresp[1:0])
    ,.bvalid(slv0_bvalid)
    ,.rid(slv0_rid[(IDWID - 1):0])
    ,.rlast(slv0_rlast)
    ,.rready(slv0_rready)
    ,.rresp(slv0_rresp[1:0])
    ,.rvalid(slv0_rvalid)
    ,.rdata(slv0_rdata[(DWID - 1):0])
    ,.wdata(slv0_wdata[(DWID - 1):0])
    ,.wlast(slv0_wlast)
    ,.wready(slv0_wready)
    ,.wstrb(slv0_wstrb[(WSTRB - 1):0])
    ,.wvalid(slv0_wvalid)


    ,.a_araddr(split102_merge200_araddr[31:0])
    ,.a_arburst(split102_merge200_arburst[1:0])
    ,.a_arextras(split102_merge200_arextras[(EXTRAS - 1):0])
    ,.a_arid(split102_merge200_arid[(IDWID - 1):0])
    ,.a_arlen(split102_merge200_arlen[7:0])
    ,.a_arready(split102_merge200_arready)
    ,.a_arvalid(split102_merge200_arvalid)
    ,.a_awaddr(split102_merge200_awaddr[31:0])
    ,.a_awburst(split102_merge200_awburst[1:0])
    ,.a_awextras(split102_merge200_awextras[(EXTRAS - 1):0])
    ,.a_awid(split102_merge200_awid[(IDWID - 1):0])
    ,.a_awlen(split102_merge200_awlen[7:0])
    ,.a_awready(split102_merge200_awready)
    ,.a_awvalid(split102_merge200_awvalid)
    ,.a_bid(split102_merge200_bid[(IDWID - 1):0])
    ,.a_bready(split102_merge200_bready)
    ,.a_bresp(split102_merge200_bresp[1:0])
    ,.a_bvalid(split102_merge200_bvalid)
    ,.a_rdata(split102_merge200_rdata[(DWID - 1):0])
    ,.a_rid(split102_merge200_rid[(IDWID - 1):0])
    ,.a_rlast(split102_merge200_rlast)
    ,.a_rready(split102_merge200_rready)
    ,.a_rresp(split102_merge200_rresp[1:0])
    ,.a_rvalid(split102_merge200_rvalid)
    ,.a_wdata(split102_merge200_wdata[(DWID - 1):0])
    ,.a_wlast(split102_merge200_wlast)
    ,.a_wready(split102_merge200_wready)
    ,.a_wstrb(split102_merge200_wstrb[(WSTRB - 1):0])
    ,.a_wvalid(split102_merge200_wvalid)

    ,.b_araddr(split103_merge200_araddr[31:0])
    ,.b_arburst(split103_merge200_arburst[1:0])
    ,.b_arextras(split103_merge200_arextras[(EXTRAS - 1):0])
    ,.b_arid(split103_merge200_arid[(IDWID - 1):0])
    ,.b_arlen(split103_merge200_arlen[7:0])
    ,.b_arready(split103_merge200_arready)
    ,.b_arvalid(split103_merge200_arvalid)
    ,.b_awaddr(split103_merge200_awaddr[31:0])
    ,.b_awburst(split103_merge200_awburst[1:0])
    ,.b_awextras(split103_merge200_awextras[(EXTRAS - 1):0])
    ,.b_awid(split103_merge200_awid[(IDWID - 1):0])
    ,.b_awlen(split103_merge200_awlen[7:0])
    ,.b_awready(split103_merge200_awready)
    ,.b_awvalid(split103_merge200_awvalid)
    ,.b_bid(split103_merge200_bid[(IDWID - 1):0])
    ,.b_bready(split103_merge200_bready)
    ,.b_bresp(split103_merge200_bresp[1:0])
    ,.b_bvalid(split103_merge200_bvalid)
    ,.b_rdata(split103_merge200_rdata[(DWID - 1):0])
    ,.b_rid(split103_merge200_rid[(IDWID - 1):0])
    ,.b_rlast(split103_merge200_rlast)
    ,.b_rready(split103_merge200_rready)
    ,.b_rresp(split103_merge200_rresp[1:0])
    ,.b_rvalid(split103_merge200_rvalid)
    ,.b_wdata(split103_merge200_wdata[(DWID - 1):0])
    ,.b_wlast(split103_merge200_wlast)
    ,.b_wready(split103_merge200_wready)
    ,.b_wstrb(split103_merge200_wstrb[(WSTRB - 1):0])
    ,.b_wvalid(split103_merge200_wvalid)

    ,.c_araddr(split108_merge200_araddr[31:0])
    ,.c_arburst(split108_merge200_arburst[1:0])
    ,.c_arextras(split108_merge200_arextras[(EXTRAS - 1):0])
    ,.c_arid(split108_merge200_arid[(IDWID - 1):0])
    ,.c_arlen(split108_merge200_arlen[7:0])
    ,.c_arready(split108_merge200_arready)
    ,.c_arvalid(split108_merge200_arvalid)
    ,.c_awaddr(split108_merge200_awaddr[31:0])
    ,.c_awburst(split108_merge200_awburst[1:0])
    ,.c_awextras(split108_merge200_awextras[(EXTRAS - 1):0])
    ,.c_awid(split108_merge200_awid[(IDWID - 1):0])
    ,.c_awlen(split108_merge200_awlen[7:0])
    ,.c_awready(split108_merge200_awready)
    ,.c_awvalid(split108_merge200_awvalid)
    ,.c_bid(split108_merge200_bid[(IDWID - 1):0])
    ,.c_bready(split108_merge200_bready)
    ,.c_bresp(split108_merge200_bresp[1:0])
    ,.c_bvalid(split108_merge200_bvalid)
    ,.c_rdata(split108_merge200_rdata[(DWID - 1):0])
    ,.c_rid(split108_merge200_rid[(IDWID - 1):0])
    ,.c_rlast(split108_merge200_rlast)
    ,.c_rready(split108_merge200_rready)
    ,.c_rresp(split108_merge200_rresp[1:0])
    ,.c_rvalid(split108_merge200_rvalid)
    ,.c_wdata(split108_merge200_wdata[(DWID - 1):0])
    ,.c_wlast(split108_merge200_wlast)
    ,.c_wready(split108_merge200_wready)
    ,.c_wstrb(split108_merge200_wstrb[(WSTRB - 1):0])
    ,.c_wvalid(split108_merge200_wvalid)

    ,.d_araddr(split111_merge200_araddr[31:0])
    ,.d_arburst(split111_merge200_arburst[1:0])
    ,.d_arextras(split111_merge200_arextras[(EXTRAS - 1):0])
    ,.d_arid(split111_merge200_arid[(IDWID - 1):0])
    ,.d_arlen(split111_merge200_arlen[7:0])
    ,.d_arready(split111_merge200_arready)
    ,.d_arvalid(split111_merge200_arvalid)
    ,.d_awaddr(split111_merge200_awaddr[31:0])
    ,.d_awburst(split111_merge200_awburst[1:0])
    ,.d_awextras(split111_merge200_awextras[(EXTRAS - 1):0])
    ,.d_awid(split111_merge200_awid[(IDWID - 1):0])
    ,.d_awlen(split111_merge200_awlen[7:0])
    ,.d_awready(split111_merge200_awready)
    ,.d_awvalid(split111_merge200_awvalid)
    ,.d_bid(split111_merge200_bid[(IDWID - 1):0])
    ,.d_bready(split111_merge200_bready)
    ,.d_bresp(split111_merge200_bresp[1:0])
    ,.d_bvalid(split111_merge200_bvalid)
    ,.d_rdata(split111_merge200_rdata[(DWID - 1):0])
    ,.d_rid(split111_merge200_rid[(IDWID - 1):0])
    ,.d_rlast(split111_merge200_rlast)
    ,.d_rready(split111_merge200_rready)
    ,.d_rresp(split111_merge200_rresp[1:0])
    ,.d_rvalid(split111_merge200_rvalid)
    ,.d_wdata(split111_merge200_wdata[(DWID - 1):0])
    ,.d_wlast(split111_merge200_wlast)
    ,.d_wready(split111_merge200_wready)
    ,.d_wstrb(split111_merge200_wstrb[(WSTRB - 1):0])
    ,.d_wvalid(split111_merge200_wvalid)
);


axi_4_merger merge207 (
     .clk(clk),.rst_n(rst_n)
    ,.araddr(slv7_araddr[31:0])
    ,.arburst(slv7_arburst[1:0])
    ,.arextras(slv7_arextras[(EXTRAS - 1):0])
    ,.arid(slv7_arid[(IDWID - 1):0])
    ,.arlen(slv7_arlen[7:0])
    ,.arready(slv7_arready)
    ,.arvalid(slv7_arvalid)
    ,.awaddr(slv7_awaddr[31:0])
    ,.awburst(slv7_awburst[1:0])
    ,.awextras(slv7_awextras[(EXTRAS - 1):0])
    ,.awid(slv7_awid[3:0])
    ,.awlen(slv7_awlen[7:0])
    ,.awready(slv7_awready)
    ,.awvalid(slv7_awvalid)
    ,.bid(slv7_bid[(IDWID - 1):0])
    ,.bready(slv7_bready)
    ,.bresp(slv7_bresp[1:0])
    ,.bvalid(slv7_bvalid)
    ,.rid(slv7_rid[(IDWID - 1):0])
    ,.rlast(slv7_rlast)
    ,.rready(slv7_rready)
    ,.rresp(slv7_rresp[1:0])
    ,.rvalid(slv7_rvalid)
    ,.rdata(slv7_rdata[(DWID - 1):0])
    ,.wdata(slv7_wdata[(DWID - 1):0])
    ,.wlast(slv7_wlast)
    ,.wready(slv7_wready)
    ,.wstrb(slv7_wstrb[(WSTRB - 1):0])
    ,.wvalid(slv7_wvalid)


    ,.a_araddr(split102_merge207_araddr[31:0])
    ,.a_arburst(split102_merge207_arburst[1:0])
    ,.a_arextras(split102_merge207_arextras[(EXTRAS - 1):0])
    ,.a_arid(split102_merge207_arid[(IDWID - 1):0])
    ,.a_arlen(split102_merge207_arlen[7:0])
    ,.a_arready(split102_merge207_arready)
    ,.a_arvalid(split102_merge207_arvalid)
    ,.a_awaddr(split102_merge207_awaddr[31:0])
    ,.a_awburst(split102_merge207_awburst[1:0])
    ,.a_awextras(split102_merge207_awextras[(EXTRAS - 1):0])
    ,.a_awid(split102_merge207_awid[(IDWID - 1):0])
    ,.a_awlen(split102_merge207_awlen[7:0])
    ,.a_awready(split102_merge207_awready)
    ,.a_awvalid(split102_merge207_awvalid)
    ,.a_bid(split102_merge207_bid[(IDWID - 1):0])
    ,.a_bready(split102_merge207_bready)
    ,.a_bresp(split102_merge207_bresp[1:0])
    ,.a_bvalid(split102_merge207_bvalid)
    ,.a_rdata(split102_merge207_rdata[(DWID - 1):0])
    ,.a_rid(split102_merge207_rid[(IDWID - 1):0])
    ,.a_rlast(split102_merge207_rlast)
    ,.a_rready(split102_merge207_rready)
    ,.a_rresp(split102_merge207_rresp[1:0])
    ,.a_rvalid(split102_merge207_rvalid)
    ,.a_wdata(split102_merge207_wdata[(DWID - 1):0])
    ,.a_wlast(split102_merge207_wlast)
    ,.a_wready(split102_merge207_wready)
    ,.a_wstrb(split102_merge207_wstrb[(WSTRB - 1):0])
    ,.a_wvalid(split102_merge207_wvalid)

    ,.b_araddr(split103_merge207_araddr[31:0])
    ,.b_arburst(split103_merge207_arburst[1:0])
    ,.b_arextras(split103_merge207_arextras[(EXTRAS - 1):0])
    ,.b_arid(split103_merge207_arid[(IDWID - 1):0])
    ,.b_arlen(split103_merge207_arlen[7:0])
    ,.b_arready(split103_merge207_arready)
    ,.b_arvalid(split103_merge207_arvalid)
    ,.b_awaddr(split103_merge207_awaddr[31:0])
    ,.b_awburst(split103_merge207_awburst[1:0])
    ,.b_awextras(split103_merge207_awextras[(EXTRAS - 1):0])
    ,.b_awid(split103_merge207_awid[(IDWID - 1):0])
    ,.b_awlen(split103_merge207_awlen[7:0])
    ,.b_awready(split103_merge207_awready)
    ,.b_awvalid(split103_merge207_awvalid)
    ,.b_bid(split103_merge207_bid[(IDWID - 1):0])
    ,.b_bready(split103_merge207_bready)
    ,.b_bresp(split103_merge207_bresp[1:0])
    ,.b_bvalid(split103_merge207_bvalid)
    ,.b_rdata(split103_merge207_rdata[(DWID - 1):0])
    ,.b_rid(split103_merge207_rid[(IDWID - 1):0])
    ,.b_rlast(split103_merge207_rlast)
    ,.b_rready(split103_merge207_rready)
    ,.b_rresp(split103_merge207_rresp[1:0])
    ,.b_rvalid(split103_merge207_rvalid)
    ,.b_wdata(split103_merge207_wdata[(DWID - 1):0])
    ,.b_wlast(split103_merge207_wlast)
    ,.b_wready(split103_merge207_wready)
    ,.b_wstrb(split103_merge207_wstrb[(WSTRB - 1):0])
    ,.b_wvalid(split103_merge207_wvalid)

    ,.c_araddr(split107_merge207_araddr[31:0])
    ,.c_arburst(split107_merge207_arburst[1:0])
    ,.c_arextras(split107_merge207_arextras[(EXTRAS - 1):0])
    ,.c_arid(split107_merge207_arid[(IDWID - 1):0])
    ,.c_arlen(split107_merge207_arlen[7:0])
    ,.c_arready(split107_merge207_arready)
    ,.c_arvalid(split107_merge207_arvalid)
    ,.c_awaddr(split107_merge207_awaddr[31:0])
    ,.c_awburst(split107_merge207_awburst[1:0])
    ,.c_awextras(split107_merge207_awextras[(EXTRAS - 1):0])
    ,.c_awid(split107_merge207_awid[(IDWID - 1):0])
    ,.c_awlen(split107_merge207_awlen[7:0])
    ,.c_awready(split107_merge207_awready)
    ,.c_awvalid(split107_merge207_awvalid)
    ,.c_bid(split107_merge207_bid[(IDWID - 1):0])
    ,.c_bready(split107_merge207_bready)
    ,.c_bresp(split107_merge207_bresp[1:0])
    ,.c_bvalid(split107_merge207_bvalid)
    ,.c_rdata(split107_merge207_rdata[(DWID - 1):0])
    ,.c_rid(split107_merge207_rid[(IDWID - 1):0])
    ,.c_rlast(split107_merge207_rlast)
    ,.c_rready(split107_merge207_rready)
    ,.c_rresp(split107_merge207_rresp[1:0])
    ,.c_rvalid(split107_merge207_rvalid)
    ,.c_wdata(split107_merge207_wdata[(DWID - 1):0])
    ,.c_wlast(split107_merge207_wlast)
    ,.c_wready(split107_merge207_wready)
    ,.c_wstrb(split107_merge207_wstrb[(WSTRB - 1):0])
    ,.c_wvalid(split107_merge207_wvalid)

    ,.d_araddr(split115_merge207_araddr[31:0])
    ,.d_arburst(split115_merge207_arburst[1:0])
    ,.d_arextras(split115_merge207_arextras[(EXTRAS - 1):0])
    ,.d_arid(split115_merge207_arid[(IDWID - 1):0])
    ,.d_arlen(split115_merge207_arlen[7:0])
    ,.d_arready(split115_merge207_arready)
    ,.d_arvalid(split115_merge207_arvalid)
    ,.d_awaddr(split115_merge207_awaddr[31:0])
    ,.d_awburst(split115_merge207_awburst[1:0])
    ,.d_awextras(split115_merge207_awextras[(EXTRAS - 1):0])
    ,.d_awid(split115_merge207_awid[(IDWID - 1):0])
    ,.d_awlen(split115_merge207_awlen[7:0])
    ,.d_awready(split115_merge207_awready)
    ,.d_awvalid(split115_merge207_awvalid)
    ,.d_bid(split115_merge207_bid[(IDWID - 1):0])
    ,.d_bready(split115_merge207_bready)
    ,.d_bresp(split115_merge207_bresp[1:0])
    ,.d_bvalid(split115_merge207_bvalid)
    ,.d_rdata(split115_merge207_rdata[(DWID - 1):0])
    ,.d_rid(split115_merge207_rid[(IDWID - 1):0])
    ,.d_rlast(split115_merge207_rlast)
    ,.d_rready(split115_merge207_rready)
    ,.d_rresp(split115_merge207_rresp[1:0])
    ,.d_rvalid(split115_merge207_rvalid)
    ,.d_wdata(split115_merge207_wdata[(DWID - 1):0])
    ,.d_wlast(split115_merge207_wlast)
    ,.d_wready(split115_merge207_wready)
    ,.d_wstrb(split115_merge207_wstrb[(WSTRB - 1):0])
    ,.d_wvalid(split115_merge207_wvalid)
);


axi_4_merger merge205 (
     .clk(clk),.rst_n(rst_n)
    ,.araddr(slv5_araddr[31:0])
    ,.arburst(slv5_arburst[1:0])
    ,.arextras(slv5_arextras[(EXTRAS - 1):0])
    ,.arid(slv5_arid[(IDWID - 1):0])
    ,.arlen(slv5_arlen[7:0])
    ,.arready(slv5_arready)
    ,.arvalid(slv5_arvalid)
    ,.awaddr(slv5_awaddr[31:0])
    ,.awburst(slv5_awburst[1:0])
    ,.awextras(slv5_awextras[(EXTRAS - 1):0])
    ,.awid(slv5_awid[3:0])
    ,.awlen(slv5_awlen[7:0])
    ,.awready(slv5_awready)
    ,.awvalid(slv5_awvalid)
    ,.bid(slv5_bid[(IDWID - 1):0])
    ,.bready(slv5_bready)
    ,.bresp(slv5_bresp[1:0])
    ,.bvalid(slv5_bvalid)
    ,.rid(slv5_rid[(IDWID - 1):0])
    ,.rlast(slv5_rlast)
    ,.rready(slv5_rready)
    ,.rresp(slv5_rresp[1:0])
    ,.rvalid(slv5_rvalid)
    ,.rdata(slv5_rdata[(DWID - 1):0])
    ,.wdata(slv5_wdata[(DWID - 1):0])
    ,.wlast(slv5_wlast)
    ,.wready(slv5_wready)
    ,.wstrb(slv5_wstrb[(WSTRB - 1):0])
    ,.wvalid(slv5_wvalid)


    ,.a_araddr(split102_merge205_araddr[31:0])
    ,.a_arburst(split102_merge205_arburst[1:0])
    ,.a_arextras(split102_merge205_arextras[(EXTRAS - 1):0])
    ,.a_arid(split102_merge205_arid[(IDWID - 1):0])
    ,.a_arlen(split102_merge205_arlen[7:0])
    ,.a_arready(split102_merge205_arready)
    ,.a_arvalid(split102_merge205_arvalid)
    ,.a_awaddr(split102_merge205_awaddr[31:0])
    ,.a_awburst(split102_merge205_awburst[1:0])
    ,.a_awextras(split102_merge205_awextras[(EXTRAS - 1):0])
    ,.a_awid(split102_merge205_awid[(IDWID - 1):0])
    ,.a_awlen(split102_merge205_awlen[7:0])
    ,.a_awready(split102_merge205_awready)
    ,.a_awvalid(split102_merge205_awvalid)
    ,.a_bid(split102_merge205_bid[(IDWID - 1):0])
    ,.a_bready(split102_merge205_bready)
    ,.a_bresp(split102_merge205_bresp[1:0])
    ,.a_bvalid(split102_merge205_bvalid)
    ,.a_rdata(split102_merge205_rdata[(DWID - 1):0])
    ,.a_rid(split102_merge205_rid[(IDWID - 1):0])
    ,.a_rlast(split102_merge205_rlast)
    ,.a_rready(split102_merge205_rready)
    ,.a_rresp(split102_merge205_rresp[1:0])
    ,.a_rvalid(split102_merge205_rvalid)
    ,.a_wdata(split102_merge205_wdata[(DWID - 1):0])
    ,.a_wlast(split102_merge205_wlast)
    ,.a_wready(split102_merge205_wready)
    ,.a_wstrb(split102_merge205_wstrb[(WSTRB - 1):0])
    ,.a_wvalid(split102_merge205_wvalid)

    ,.b_araddr(split106_merge205_araddr[31:0])
    ,.b_arburst(split106_merge205_arburst[1:0])
    ,.b_arextras(split106_merge205_arextras[(EXTRAS - 1):0])
    ,.b_arid(split106_merge205_arid[(IDWID - 1):0])
    ,.b_arlen(split106_merge205_arlen[7:0])
    ,.b_arready(split106_merge205_arready)
    ,.b_arvalid(split106_merge205_arvalid)
    ,.b_awaddr(split106_merge205_awaddr[31:0])
    ,.b_awburst(split106_merge205_awburst[1:0])
    ,.b_awextras(split106_merge205_awextras[(EXTRAS - 1):0])
    ,.b_awid(split106_merge205_awid[(IDWID - 1):0])
    ,.b_awlen(split106_merge205_awlen[7:0])
    ,.b_awready(split106_merge205_awready)
    ,.b_awvalid(split106_merge205_awvalid)
    ,.b_bid(split106_merge205_bid[(IDWID - 1):0])
    ,.b_bready(split106_merge205_bready)
    ,.b_bresp(split106_merge205_bresp[1:0])
    ,.b_bvalid(split106_merge205_bvalid)
    ,.b_rdata(split106_merge205_rdata[(DWID - 1):0])
    ,.b_rid(split106_merge205_rid[(IDWID - 1):0])
    ,.b_rlast(split106_merge205_rlast)
    ,.b_rready(split106_merge205_rready)
    ,.b_rresp(split106_merge205_rresp[1:0])
    ,.b_rvalid(split106_merge205_rvalid)
    ,.b_wdata(split106_merge205_wdata[(DWID - 1):0])
    ,.b_wlast(split106_merge205_wlast)
    ,.b_wready(split106_merge205_wready)
    ,.b_wstrb(split106_merge205_wstrb[(WSTRB - 1):0])
    ,.b_wvalid(split106_merge205_wvalid)

    ,.c_araddr(split108_merge205_araddr[31:0])
    ,.c_arburst(split108_merge205_arburst[1:0])
    ,.c_arextras(split108_merge205_arextras[(EXTRAS - 1):0])
    ,.c_arid(split108_merge205_arid[(IDWID - 1):0])
    ,.c_arlen(split108_merge205_arlen[7:0])
    ,.c_arready(split108_merge205_arready)
    ,.c_arvalid(split108_merge205_arvalid)
    ,.c_awaddr(split108_merge205_awaddr[31:0])
    ,.c_awburst(split108_merge205_awburst[1:0])
    ,.c_awextras(split108_merge205_awextras[(EXTRAS - 1):0])
    ,.c_awid(split108_merge205_awid[(IDWID - 1):0])
    ,.c_awlen(split108_merge205_awlen[7:0])
    ,.c_awready(split108_merge205_awready)
    ,.c_awvalid(split108_merge205_awvalid)
    ,.c_bid(split108_merge205_bid[(IDWID - 1):0])
    ,.c_bready(split108_merge205_bready)
    ,.c_bresp(split108_merge205_bresp[1:0])
    ,.c_bvalid(split108_merge205_bvalid)
    ,.c_rdata(split108_merge205_rdata[(DWID - 1):0])
    ,.c_rid(split108_merge205_rid[(IDWID - 1):0])
    ,.c_rlast(split108_merge205_rlast)
    ,.c_rready(split108_merge205_rready)
    ,.c_rresp(split108_merge205_rresp[1:0])
    ,.c_rvalid(split108_merge205_rvalid)
    ,.c_wdata(split108_merge205_wdata[(DWID - 1):0])
    ,.c_wlast(split108_merge205_wlast)
    ,.c_wready(split108_merge205_wready)
    ,.c_wstrb(split108_merge205_wstrb[(WSTRB - 1):0])
    ,.c_wvalid(split108_merge205_wvalid)

    ,.d_araddr(split113_merge205_araddr[31:0])
    ,.d_arburst(split113_merge205_arburst[1:0])
    ,.d_arextras(split113_merge205_arextras[(EXTRAS - 1):0])
    ,.d_arid(split113_merge205_arid[(IDWID - 1):0])
    ,.d_arlen(split113_merge205_arlen[7:0])
    ,.d_arready(split113_merge205_arready)
    ,.d_arvalid(split113_merge205_arvalid)
    ,.d_awaddr(split113_merge205_awaddr[31:0])
    ,.d_awburst(split113_merge205_awburst[1:0])
    ,.d_awextras(split113_merge205_awextras[(EXTRAS - 1):0])
    ,.d_awid(split113_merge205_awid[(IDWID - 1):0])
    ,.d_awlen(split113_merge205_awlen[7:0])
    ,.d_awready(split113_merge205_awready)
    ,.d_awvalid(split113_merge205_awvalid)
    ,.d_bid(split113_merge205_bid[(IDWID - 1):0])
    ,.d_bready(split113_merge205_bready)
    ,.d_bresp(split113_merge205_bresp[1:0])
    ,.d_bvalid(split113_merge205_bvalid)
    ,.d_rdata(split113_merge205_rdata[(DWID - 1):0])
    ,.d_rid(split113_merge205_rid[(IDWID - 1):0])
    ,.d_rlast(split113_merge205_rlast)
    ,.d_rready(split113_merge205_rready)
    ,.d_rresp(split113_merge205_rresp[1:0])
    ,.d_rvalid(split113_merge205_rvalid)
    ,.d_wdata(split113_merge205_wdata[(DWID - 1):0])
    ,.d_wlast(split113_merge205_wlast)
    ,.d_wready(split113_merge205_wready)
    ,.d_wstrb(split113_merge205_wstrb[(WSTRB - 1):0])
    ,.d_wvalid(split113_merge205_wvalid)
);


axi_4_merger merge213 (
     .clk(clk),.rst_n(rst_n)
    ,.araddr(slv13_araddr[31:0])
    ,.arburst(slv13_arburst[1:0])
    ,.arextras(slv13_arextras[(EXTRAS - 1):0])
    ,.arid(slv13_arid[(IDWID - 1):0])
    ,.arlen(slv13_arlen[7:0])
    ,.arready(slv13_arready)
    ,.arvalid(slv13_arvalid)
    ,.awaddr(slv13_awaddr[31:0])
    ,.awburst(slv13_awburst[1:0])
    ,.awextras(slv13_awextras[(EXTRAS - 1):0])
    ,.awid(slv13_awid[3:0])
    ,.awlen(slv13_awlen[7:0])
    ,.awready(slv13_awready)
    ,.awvalid(slv13_awvalid)
    ,.bid(slv13_bid[(IDWID - 1):0])
    ,.bready(slv13_bready)
    ,.bresp(slv13_bresp[1:0])
    ,.bvalid(slv13_bvalid)
    ,.rid(slv13_rid[(IDWID - 1):0])
    ,.rlast(slv13_rlast)
    ,.rready(slv13_rready)
    ,.rresp(slv13_rresp[1:0])
    ,.rvalid(slv13_rvalid)
    ,.rdata(slv13_rdata[(DWID - 1):0])
    ,.wdata(slv13_wdata[(DWID - 1):0])
    ,.wlast(slv13_wlast)
    ,.wready(slv13_wready)
    ,.wstrb(slv13_wstrb[(WSTRB - 1):0])
    ,.wvalid(slv13_wvalid)


    ,.a_araddr(split104_merge213_araddr[31:0])
    ,.a_arburst(split104_merge213_arburst[1:0])
    ,.a_arextras(split104_merge213_arextras[(EXTRAS - 1):0])
    ,.a_arid(split104_merge213_arid[(IDWID - 1):0])
    ,.a_arlen(split104_merge213_arlen[7:0])
    ,.a_arready(split104_merge213_arready)
    ,.a_arvalid(split104_merge213_arvalid)
    ,.a_awaddr(split104_merge213_awaddr[31:0])
    ,.a_awburst(split104_merge213_awburst[1:0])
    ,.a_awextras(split104_merge213_awextras[(EXTRAS - 1):0])
    ,.a_awid(split104_merge213_awid[(IDWID - 1):0])
    ,.a_awlen(split104_merge213_awlen[7:0])
    ,.a_awready(split104_merge213_awready)
    ,.a_awvalid(split104_merge213_awvalid)
    ,.a_bid(split104_merge213_bid[(IDWID - 1):0])
    ,.a_bready(split104_merge213_bready)
    ,.a_bresp(split104_merge213_bresp[1:0])
    ,.a_bvalid(split104_merge213_bvalid)
    ,.a_rdata(split104_merge213_rdata[(DWID - 1):0])
    ,.a_rid(split104_merge213_rid[(IDWID - 1):0])
    ,.a_rlast(split104_merge213_rlast)
    ,.a_rready(split104_merge213_rready)
    ,.a_rresp(split104_merge213_rresp[1:0])
    ,.a_rvalid(split104_merge213_rvalid)
    ,.a_wdata(split104_merge213_wdata[(DWID - 1):0])
    ,.a_wlast(split104_merge213_wlast)
    ,.a_wready(split104_merge213_wready)
    ,.a_wstrb(split104_merge213_wstrb[(WSTRB - 1):0])
    ,.a_wvalid(split104_merge213_wvalid)

    ,.b_araddr(split105_merge213_araddr[31:0])
    ,.b_arburst(split105_merge213_arburst[1:0])
    ,.b_arextras(split105_merge213_arextras[(EXTRAS - 1):0])
    ,.b_arid(split105_merge213_arid[(IDWID - 1):0])
    ,.b_arlen(split105_merge213_arlen[7:0])
    ,.b_arready(split105_merge213_arready)
    ,.b_arvalid(split105_merge213_arvalid)
    ,.b_awaddr(split105_merge213_awaddr[31:0])
    ,.b_awburst(split105_merge213_awburst[1:0])
    ,.b_awextras(split105_merge213_awextras[(EXTRAS - 1):0])
    ,.b_awid(split105_merge213_awid[(IDWID - 1):0])
    ,.b_awlen(split105_merge213_awlen[7:0])
    ,.b_awready(split105_merge213_awready)
    ,.b_awvalid(split105_merge213_awvalid)
    ,.b_bid(split105_merge213_bid[(IDWID - 1):0])
    ,.b_bready(split105_merge213_bready)
    ,.b_bresp(split105_merge213_bresp[1:0])
    ,.b_bvalid(split105_merge213_bvalid)
    ,.b_rdata(split105_merge213_rdata[(DWID - 1):0])
    ,.b_rid(split105_merge213_rid[(IDWID - 1):0])
    ,.b_rlast(split105_merge213_rlast)
    ,.b_rready(split105_merge213_rready)
    ,.b_rresp(split105_merge213_rresp[1:0])
    ,.b_rvalid(split105_merge213_rvalid)
    ,.b_wdata(split105_merge213_wdata[(DWID - 1):0])
    ,.b_wlast(split105_merge213_wlast)
    ,.b_wready(split105_merge213_wready)
    ,.b_wstrb(split105_merge213_wstrb[(WSTRB - 1):0])
    ,.b_wvalid(split105_merge213_wvalid)

    ,.c_araddr(split106_merge213_araddr[31:0])
    ,.c_arburst(split106_merge213_arburst[1:0])
    ,.c_arextras(split106_merge213_arextras[(EXTRAS - 1):0])
    ,.c_arid(split106_merge213_arid[(IDWID - 1):0])
    ,.c_arlen(split106_merge213_arlen[7:0])
    ,.c_arready(split106_merge213_arready)
    ,.c_arvalid(split106_merge213_arvalid)
    ,.c_awaddr(split106_merge213_awaddr[31:0])
    ,.c_awburst(split106_merge213_awburst[1:0])
    ,.c_awextras(split106_merge213_awextras[(EXTRAS - 1):0])
    ,.c_awid(split106_merge213_awid[(IDWID - 1):0])
    ,.c_awlen(split106_merge213_awlen[7:0])
    ,.c_awready(split106_merge213_awready)
    ,.c_awvalid(split106_merge213_awvalid)
    ,.c_bid(split106_merge213_bid[(IDWID - 1):0])
    ,.c_bready(split106_merge213_bready)
    ,.c_bresp(split106_merge213_bresp[1:0])
    ,.c_bvalid(split106_merge213_bvalid)
    ,.c_rdata(split106_merge213_rdata[(DWID - 1):0])
    ,.c_rid(split106_merge213_rid[(IDWID - 1):0])
    ,.c_rlast(split106_merge213_rlast)
    ,.c_rready(split106_merge213_rready)
    ,.c_rresp(split106_merge213_rresp[1:0])
    ,.c_rvalid(split106_merge213_rvalid)
    ,.c_wdata(split106_merge213_wdata[(DWID - 1):0])
    ,.c_wlast(split106_merge213_wlast)
    ,.c_wready(split106_merge213_wready)
    ,.c_wstrb(split106_merge213_wstrb[(WSTRB - 1):0])
    ,.c_wvalid(split106_merge213_wvalid)

    ,.d_araddr(split111_merge213_araddr[31:0])
    ,.d_arburst(split111_merge213_arburst[1:0])
    ,.d_arextras(split111_merge213_arextras[(EXTRAS - 1):0])
    ,.d_arid(split111_merge213_arid[(IDWID - 1):0])
    ,.d_arlen(split111_merge213_arlen[7:0])
    ,.d_arready(split111_merge213_arready)
    ,.d_arvalid(split111_merge213_arvalid)
    ,.d_awaddr(split111_merge213_awaddr[31:0])
    ,.d_awburst(split111_merge213_awburst[1:0])
    ,.d_awextras(split111_merge213_awextras[(EXTRAS - 1):0])
    ,.d_awid(split111_merge213_awid[(IDWID - 1):0])
    ,.d_awlen(split111_merge213_awlen[7:0])
    ,.d_awready(split111_merge213_awready)
    ,.d_awvalid(split111_merge213_awvalid)
    ,.d_bid(split111_merge213_bid[(IDWID - 1):0])
    ,.d_bready(split111_merge213_bready)
    ,.d_bresp(split111_merge213_bresp[1:0])
    ,.d_bvalid(split111_merge213_bvalid)
    ,.d_rdata(split111_merge213_rdata[(DWID - 1):0])
    ,.d_rid(split111_merge213_rid[(IDWID - 1):0])
    ,.d_rlast(split111_merge213_rlast)
    ,.d_rready(split111_merge213_rready)
    ,.d_rresp(split111_merge213_rresp[1:0])
    ,.d_rvalid(split111_merge213_rvalid)
    ,.d_wdata(split111_merge213_wdata[(DWID - 1):0])
    ,.d_wlast(split111_merge213_wlast)
    ,.d_wready(split111_merge213_wready)
    ,.d_wstrb(split111_merge213_wstrb[(WSTRB - 1):0])
    ,.d_wvalid(split111_merge213_wvalid)
);


axi_4_merger merge214 (
     .clk(clk),.rst_n(rst_n)
    ,.araddr(slv14_araddr[31:0])
    ,.arburst(slv14_arburst[1:0])
    ,.arextras(slv14_arextras[(EXTRAS - 1):0])
    ,.arid(slv14_arid[(IDWID - 1):0])
    ,.arlen(slv14_arlen[7:0])
    ,.arready(slv14_arready)
    ,.arvalid(slv14_arvalid)
    ,.awaddr(slv14_awaddr[31:0])
    ,.awburst(slv14_awburst[1:0])
    ,.awextras(slv14_awextras[(EXTRAS - 1):0])
    ,.awid(slv14_awid[3:0])
    ,.awlen(slv14_awlen[7:0])
    ,.awready(slv14_awready)
    ,.awvalid(slv14_awvalid)
    ,.bid(slv14_bid[(IDWID - 1):0])
    ,.bready(slv14_bready)
    ,.bresp(slv14_bresp[1:0])
    ,.bvalid(slv14_bvalid)
    ,.rid(slv14_rid[(IDWID - 1):0])
    ,.rlast(slv14_rlast)
    ,.rready(slv14_rready)
    ,.rresp(slv14_rresp[1:0])
    ,.rvalid(slv14_rvalid)
    ,.rdata(slv14_rdata[(DWID - 1):0])
    ,.wdata(slv14_wdata[(DWID - 1):0])
    ,.wlast(slv14_wlast)
    ,.wready(slv14_wready)
    ,.wstrb(slv14_wstrb[(WSTRB - 1):0])
    ,.wvalid(slv14_wvalid)


    ,.a_araddr(split104_merge214_araddr[31:0])
    ,.a_arburst(split104_merge214_arburst[1:0])
    ,.a_arextras(split104_merge214_arextras[(EXTRAS - 1):0])
    ,.a_arid(split104_merge214_arid[(IDWID - 1):0])
    ,.a_arlen(split104_merge214_arlen[7:0])
    ,.a_arready(split104_merge214_arready)
    ,.a_arvalid(split104_merge214_arvalid)
    ,.a_awaddr(split104_merge214_awaddr[31:0])
    ,.a_awburst(split104_merge214_awburst[1:0])
    ,.a_awextras(split104_merge214_awextras[(EXTRAS - 1):0])
    ,.a_awid(split104_merge214_awid[(IDWID - 1):0])
    ,.a_awlen(split104_merge214_awlen[7:0])
    ,.a_awready(split104_merge214_awready)
    ,.a_awvalid(split104_merge214_awvalid)
    ,.a_bid(split104_merge214_bid[(IDWID - 1):0])
    ,.a_bready(split104_merge214_bready)
    ,.a_bresp(split104_merge214_bresp[1:0])
    ,.a_bvalid(split104_merge214_bvalid)
    ,.a_rdata(split104_merge214_rdata[(DWID - 1):0])
    ,.a_rid(split104_merge214_rid[(IDWID - 1):0])
    ,.a_rlast(split104_merge214_rlast)
    ,.a_rready(split104_merge214_rready)
    ,.a_rresp(split104_merge214_rresp[1:0])
    ,.a_rvalid(split104_merge214_rvalid)
    ,.a_wdata(split104_merge214_wdata[(DWID - 1):0])
    ,.a_wlast(split104_merge214_wlast)
    ,.a_wready(split104_merge214_wready)
    ,.a_wstrb(split104_merge214_wstrb[(WSTRB - 1):0])
    ,.a_wvalid(split104_merge214_wvalid)

    ,.b_araddr(split110_merge214_araddr[31:0])
    ,.b_arburst(split110_merge214_arburst[1:0])
    ,.b_arextras(split110_merge214_arextras[(EXTRAS - 1):0])
    ,.b_arid(split110_merge214_arid[(IDWID - 1):0])
    ,.b_arlen(split110_merge214_arlen[7:0])
    ,.b_arready(split110_merge214_arready)
    ,.b_arvalid(split110_merge214_arvalid)
    ,.b_awaddr(split110_merge214_awaddr[31:0])
    ,.b_awburst(split110_merge214_awburst[1:0])
    ,.b_awextras(split110_merge214_awextras[(EXTRAS - 1):0])
    ,.b_awid(split110_merge214_awid[(IDWID - 1):0])
    ,.b_awlen(split110_merge214_awlen[7:0])
    ,.b_awready(split110_merge214_awready)
    ,.b_awvalid(split110_merge214_awvalid)
    ,.b_bid(split110_merge214_bid[(IDWID - 1):0])
    ,.b_bready(split110_merge214_bready)
    ,.b_bresp(split110_merge214_bresp[1:0])
    ,.b_bvalid(split110_merge214_bvalid)
    ,.b_rdata(split110_merge214_rdata[(DWID - 1):0])
    ,.b_rid(split110_merge214_rid[(IDWID - 1):0])
    ,.b_rlast(split110_merge214_rlast)
    ,.b_rready(split110_merge214_rready)
    ,.b_rresp(split110_merge214_rresp[1:0])
    ,.b_rvalid(split110_merge214_rvalid)
    ,.b_wdata(split110_merge214_wdata[(DWID - 1):0])
    ,.b_wlast(split110_merge214_wlast)
    ,.b_wready(split110_merge214_wready)
    ,.b_wstrb(split110_merge214_wstrb[(WSTRB - 1):0])
    ,.b_wvalid(split110_merge214_wvalid)

    ,.c_araddr(split111_merge214_araddr[31:0])
    ,.c_arburst(split111_merge214_arburst[1:0])
    ,.c_arextras(split111_merge214_arextras[(EXTRAS - 1):0])
    ,.c_arid(split111_merge214_arid[(IDWID - 1):0])
    ,.c_arlen(split111_merge214_arlen[7:0])
    ,.c_arready(split111_merge214_arready)
    ,.c_arvalid(split111_merge214_arvalid)
    ,.c_awaddr(split111_merge214_awaddr[31:0])
    ,.c_awburst(split111_merge214_awburst[1:0])
    ,.c_awextras(split111_merge214_awextras[(EXTRAS - 1):0])
    ,.c_awid(split111_merge214_awid[(IDWID - 1):0])
    ,.c_awlen(split111_merge214_awlen[7:0])
    ,.c_awready(split111_merge214_awready)
    ,.c_awvalid(split111_merge214_awvalid)
    ,.c_bid(split111_merge214_bid[(IDWID - 1):0])
    ,.c_bready(split111_merge214_bready)
    ,.c_bresp(split111_merge214_bresp[1:0])
    ,.c_bvalid(split111_merge214_bvalid)
    ,.c_rdata(split111_merge214_rdata[(DWID - 1):0])
    ,.c_rid(split111_merge214_rid[(IDWID - 1):0])
    ,.c_rlast(split111_merge214_rlast)
    ,.c_rready(split111_merge214_rready)
    ,.c_rresp(split111_merge214_rresp[1:0])
    ,.c_rvalid(split111_merge214_rvalid)
    ,.c_wdata(split111_merge214_wdata[(DWID - 1):0])
    ,.c_wlast(split111_merge214_wlast)
    ,.c_wready(split111_merge214_wready)
    ,.c_wstrb(split111_merge214_wstrb[(WSTRB - 1):0])
    ,.c_wvalid(split111_merge214_wvalid)

    ,.d_araddr(split115_merge214_araddr[31:0])
    ,.d_arburst(split115_merge214_arburst[1:0])
    ,.d_arextras(split115_merge214_arextras[(EXTRAS - 1):0])
    ,.d_arid(split115_merge214_arid[(IDWID - 1):0])
    ,.d_arlen(split115_merge214_arlen[7:0])
    ,.d_arready(split115_merge214_arready)
    ,.d_arvalid(split115_merge214_arvalid)
    ,.d_awaddr(split115_merge214_awaddr[31:0])
    ,.d_awburst(split115_merge214_awburst[1:0])
    ,.d_awextras(split115_merge214_awextras[(EXTRAS - 1):0])
    ,.d_awid(split115_merge214_awid[(IDWID - 1):0])
    ,.d_awlen(split115_merge214_awlen[7:0])
    ,.d_awready(split115_merge214_awready)
    ,.d_awvalid(split115_merge214_awvalid)
    ,.d_bid(split115_merge214_bid[(IDWID - 1):0])
    ,.d_bready(split115_merge214_bready)
    ,.d_bresp(split115_merge214_bresp[1:0])
    ,.d_bvalid(split115_merge214_bvalid)
    ,.d_rdata(split115_merge214_rdata[(DWID - 1):0])
    ,.d_rid(split115_merge214_rid[(IDWID - 1):0])
    ,.d_rlast(split115_merge214_rlast)
    ,.d_rready(split115_merge214_rready)
    ,.d_rresp(split115_merge214_rresp[1:0])
    ,.d_rvalid(split115_merge214_rvalid)
    ,.d_wdata(split115_merge214_wdata[(DWID - 1):0])
    ,.d_wlast(split115_merge214_wlast)
    ,.d_wready(split115_merge214_wready)
    ,.d_wstrb(split115_merge214_wstrb[(WSTRB - 1):0])
    ,.d_wvalid(split115_merge214_wvalid)
);


axi_4_merger merge204 (
     .clk(clk),.rst_n(rst_n)
    ,.araddr(slv4_araddr[31:0])
    ,.arburst(slv4_arburst[1:0])
    ,.arextras(slv4_arextras[(EXTRAS - 1):0])
    ,.arid(slv4_arid[(IDWID - 1):0])
    ,.arlen(slv4_arlen[7:0])
    ,.arready(slv4_arready)
    ,.arvalid(slv4_arvalid)
    ,.awaddr(slv4_awaddr[31:0])
    ,.awburst(slv4_awburst[1:0])
    ,.awextras(slv4_awextras[(EXTRAS - 1):0])
    ,.awid(slv4_awid[3:0])
    ,.awlen(slv4_awlen[7:0])
    ,.awready(slv4_awready)
    ,.awvalid(slv4_awvalid)
    ,.bid(slv4_bid[(IDWID - 1):0])
    ,.bready(slv4_bready)
    ,.bresp(slv4_bresp[1:0])
    ,.bvalid(slv4_bvalid)
    ,.rid(slv4_rid[(IDWID - 1):0])
    ,.rlast(slv4_rlast)
    ,.rready(slv4_rready)
    ,.rresp(slv4_rresp[1:0])
    ,.rvalid(slv4_rvalid)
    ,.rdata(slv4_rdata[(DWID - 1):0])
    ,.wdata(slv4_wdata[(DWID - 1):0])
    ,.wlast(slv4_wlast)
    ,.wready(slv4_wready)
    ,.wstrb(slv4_wstrb[(WSTRB - 1):0])
    ,.wvalid(slv4_wvalid)


    ,.a_araddr(split105_merge204_araddr[31:0])
    ,.a_arburst(split105_merge204_arburst[1:0])
    ,.a_arextras(split105_merge204_arextras[(EXTRAS - 1):0])
    ,.a_arid(split105_merge204_arid[(IDWID - 1):0])
    ,.a_arlen(split105_merge204_arlen[7:0])
    ,.a_arready(split105_merge204_arready)
    ,.a_arvalid(split105_merge204_arvalid)
    ,.a_awaddr(split105_merge204_awaddr[31:0])
    ,.a_awburst(split105_merge204_awburst[1:0])
    ,.a_awextras(split105_merge204_awextras[(EXTRAS - 1):0])
    ,.a_awid(split105_merge204_awid[(IDWID - 1):0])
    ,.a_awlen(split105_merge204_awlen[7:0])
    ,.a_awready(split105_merge204_awready)
    ,.a_awvalid(split105_merge204_awvalid)
    ,.a_bid(split105_merge204_bid[(IDWID - 1):0])
    ,.a_bready(split105_merge204_bready)
    ,.a_bresp(split105_merge204_bresp[1:0])
    ,.a_bvalid(split105_merge204_bvalid)
    ,.a_rdata(split105_merge204_rdata[(DWID - 1):0])
    ,.a_rid(split105_merge204_rid[(IDWID - 1):0])
    ,.a_rlast(split105_merge204_rlast)
    ,.a_rready(split105_merge204_rready)
    ,.a_rresp(split105_merge204_rresp[1:0])
    ,.a_rvalid(split105_merge204_rvalid)
    ,.a_wdata(split105_merge204_wdata[(DWID - 1):0])
    ,.a_wlast(split105_merge204_wlast)
    ,.a_wready(split105_merge204_wready)
    ,.a_wstrb(split105_merge204_wstrb[(WSTRB - 1):0])
    ,.a_wvalid(split105_merge204_wvalid)

    ,.b_araddr(split106_merge204_araddr[31:0])
    ,.b_arburst(split106_merge204_arburst[1:0])
    ,.b_arextras(split106_merge204_arextras[(EXTRAS - 1):0])
    ,.b_arid(split106_merge204_arid[(IDWID - 1):0])
    ,.b_arlen(split106_merge204_arlen[7:0])
    ,.b_arready(split106_merge204_arready)
    ,.b_arvalid(split106_merge204_arvalid)
    ,.b_awaddr(split106_merge204_awaddr[31:0])
    ,.b_awburst(split106_merge204_awburst[1:0])
    ,.b_awextras(split106_merge204_awextras[(EXTRAS - 1):0])
    ,.b_awid(split106_merge204_awid[(IDWID - 1):0])
    ,.b_awlen(split106_merge204_awlen[7:0])
    ,.b_awready(split106_merge204_awready)
    ,.b_awvalid(split106_merge204_awvalid)
    ,.b_bid(split106_merge204_bid[(IDWID - 1):0])
    ,.b_bready(split106_merge204_bready)
    ,.b_bresp(split106_merge204_bresp[1:0])
    ,.b_bvalid(split106_merge204_bvalid)
    ,.b_rdata(split106_merge204_rdata[(DWID - 1):0])
    ,.b_rid(split106_merge204_rid[(IDWID - 1):0])
    ,.b_rlast(split106_merge204_rlast)
    ,.b_rready(split106_merge204_rready)
    ,.b_rresp(split106_merge204_rresp[1:0])
    ,.b_rvalid(split106_merge204_rvalid)
    ,.b_wdata(split106_merge204_wdata[(DWID - 1):0])
    ,.b_wlast(split106_merge204_wlast)
    ,.b_wready(split106_merge204_wready)
    ,.b_wstrb(split106_merge204_wstrb[(WSTRB - 1):0])
    ,.b_wvalid(split106_merge204_wvalid)

    ,.c_araddr(split109_merge204_araddr[31:0])
    ,.c_arburst(split109_merge204_arburst[1:0])
    ,.c_arextras(split109_merge204_arextras[(EXTRAS - 1):0])
    ,.c_arid(split109_merge204_arid[(IDWID - 1):0])
    ,.c_arlen(split109_merge204_arlen[7:0])
    ,.c_arready(split109_merge204_arready)
    ,.c_arvalid(split109_merge204_arvalid)
    ,.c_awaddr(split109_merge204_awaddr[31:0])
    ,.c_awburst(split109_merge204_awburst[1:0])
    ,.c_awextras(split109_merge204_awextras[(EXTRAS - 1):0])
    ,.c_awid(split109_merge204_awid[(IDWID - 1):0])
    ,.c_awlen(split109_merge204_awlen[7:0])
    ,.c_awready(split109_merge204_awready)
    ,.c_awvalid(split109_merge204_awvalid)
    ,.c_bid(split109_merge204_bid[(IDWID - 1):0])
    ,.c_bready(split109_merge204_bready)
    ,.c_bresp(split109_merge204_bresp[1:0])
    ,.c_bvalid(split109_merge204_bvalid)
    ,.c_rdata(split109_merge204_rdata[(DWID - 1):0])
    ,.c_rid(split109_merge204_rid[(IDWID - 1):0])
    ,.c_rlast(split109_merge204_rlast)
    ,.c_rready(split109_merge204_rready)
    ,.c_rresp(split109_merge204_rresp[1:0])
    ,.c_rvalid(split109_merge204_rvalid)
    ,.c_wdata(split109_merge204_wdata[(DWID - 1):0])
    ,.c_wlast(split109_merge204_wlast)
    ,.c_wready(split109_merge204_wready)
    ,.c_wstrb(split109_merge204_wstrb[(WSTRB - 1):0])
    ,.c_wvalid(split109_merge204_wvalid)

    ,.d_araddr(split114_merge204_araddr[31:0])
    ,.d_arburst(split114_merge204_arburst[1:0])
    ,.d_arextras(split114_merge204_arextras[(EXTRAS - 1):0])
    ,.d_arid(split114_merge204_arid[(IDWID - 1):0])
    ,.d_arlen(split114_merge204_arlen[7:0])
    ,.d_arready(split114_merge204_arready)
    ,.d_arvalid(split114_merge204_arvalid)
    ,.d_awaddr(split114_merge204_awaddr[31:0])
    ,.d_awburst(split114_merge204_awburst[1:0])
    ,.d_awextras(split114_merge204_awextras[(EXTRAS - 1):0])
    ,.d_awid(split114_merge204_awid[(IDWID - 1):0])
    ,.d_awlen(split114_merge204_awlen[7:0])
    ,.d_awready(split114_merge204_awready)
    ,.d_awvalid(split114_merge204_awvalid)
    ,.d_bid(split114_merge204_bid[(IDWID - 1):0])
    ,.d_bready(split114_merge204_bready)
    ,.d_bresp(split114_merge204_bresp[1:0])
    ,.d_bvalid(split114_merge204_bvalid)
    ,.d_rdata(split114_merge204_rdata[(DWID - 1):0])
    ,.d_rid(split114_merge204_rid[(IDWID - 1):0])
    ,.d_rlast(split114_merge204_rlast)
    ,.d_rready(split114_merge204_rready)
    ,.d_rresp(split114_merge204_rresp[1:0])
    ,.d_rvalid(split114_merge204_rvalid)
    ,.d_wdata(split114_merge204_wdata[(DWID - 1):0])
    ,.d_wlast(split114_merge204_wlast)
    ,.d_wready(split114_merge204_wready)
    ,.d_wstrb(split114_merge204_wstrb[(WSTRB - 1):0])
    ,.d_wvalid(split114_merge204_wvalid)
);


axi_4_merger merge210 (
     .clk(clk),.rst_n(rst_n)
    ,.araddr(slv10_araddr[31:0])
    ,.arburst(slv10_arburst[1:0])
    ,.arextras(slv10_arextras[(EXTRAS - 1):0])
    ,.arid(slv10_arid[(IDWID - 1):0])
    ,.arlen(slv10_arlen[7:0])
    ,.arready(slv10_arready)
    ,.arvalid(slv10_arvalid)
    ,.awaddr(slv10_awaddr[31:0])
    ,.awburst(slv10_awburst[1:0])
    ,.awextras(slv10_awextras[(EXTRAS - 1):0])
    ,.awid(slv10_awid[3:0])
    ,.awlen(slv10_awlen[7:0])
    ,.awready(slv10_awready)
    ,.awvalid(slv10_awvalid)
    ,.bid(slv10_bid[(IDWID - 1):0])
    ,.bready(slv10_bready)
    ,.bresp(slv10_bresp[1:0])
    ,.bvalid(slv10_bvalid)
    ,.rid(slv10_rid[(IDWID - 1):0])
    ,.rlast(slv10_rlast)
    ,.rready(slv10_rready)
    ,.rresp(slv10_rresp[1:0])
    ,.rvalid(slv10_rvalid)
    ,.rdata(slv10_rdata[(DWID - 1):0])
    ,.wdata(slv10_wdata[(DWID - 1):0])
    ,.wlast(slv10_wlast)
    ,.wready(slv10_wready)
    ,.wstrb(slv10_wstrb[(WSTRB - 1):0])
    ,.wvalid(slv10_wvalid)


    ,.a_araddr(split107_merge210_araddr[31:0])
    ,.a_arburst(split107_merge210_arburst[1:0])
    ,.a_arextras(split107_merge210_arextras[(EXTRAS - 1):0])
    ,.a_arid(split107_merge210_arid[(IDWID - 1):0])
    ,.a_arlen(split107_merge210_arlen[7:0])
    ,.a_arready(split107_merge210_arready)
    ,.a_arvalid(split107_merge210_arvalid)
    ,.a_awaddr(split107_merge210_awaddr[31:0])
    ,.a_awburst(split107_merge210_awburst[1:0])
    ,.a_awextras(split107_merge210_awextras[(EXTRAS - 1):0])
    ,.a_awid(split107_merge210_awid[(IDWID - 1):0])
    ,.a_awlen(split107_merge210_awlen[7:0])
    ,.a_awready(split107_merge210_awready)
    ,.a_awvalid(split107_merge210_awvalid)
    ,.a_bid(split107_merge210_bid[(IDWID - 1):0])
    ,.a_bready(split107_merge210_bready)
    ,.a_bresp(split107_merge210_bresp[1:0])
    ,.a_bvalid(split107_merge210_bvalid)
    ,.a_rdata(split107_merge210_rdata[(DWID - 1):0])
    ,.a_rid(split107_merge210_rid[(IDWID - 1):0])
    ,.a_rlast(split107_merge210_rlast)
    ,.a_rready(split107_merge210_rready)
    ,.a_rresp(split107_merge210_rresp[1:0])
    ,.a_rvalid(split107_merge210_rvalid)
    ,.a_wdata(split107_merge210_wdata[(DWID - 1):0])
    ,.a_wlast(split107_merge210_wlast)
    ,.a_wready(split107_merge210_wready)
    ,.a_wstrb(split107_merge210_wstrb[(WSTRB - 1):0])
    ,.a_wvalid(split107_merge210_wvalid)

    ,.b_araddr(split112_merge210_araddr[31:0])
    ,.b_arburst(split112_merge210_arburst[1:0])
    ,.b_arextras(split112_merge210_arextras[(EXTRAS - 1):0])
    ,.b_arid(split112_merge210_arid[(IDWID - 1):0])
    ,.b_arlen(split112_merge210_arlen[7:0])
    ,.b_arready(split112_merge210_arready)
    ,.b_arvalid(split112_merge210_arvalid)
    ,.b_awaddr(split112_merge210_awaddr[31:0])
    ,.b_awburst(split112_merge210_awburst[1:0])
    ,.b_awextras(split112_merge210_awextras[(EXTRAS - 1):0])
    ,.b_awid(split112_merge210_awid[(IDWID - 1):0])
    ,.b_awlen(split112_merge210_awlen[7:0])
    ,.b_awready(split112_merge210_awready)
    ,.b_awvalid(split112_merge210_awvalid)
    ,.b_bid(split112_merge210_bid[(IDWID - 1):0])
    ,.b_bready(split112_merge210_bready)
    ,.b_bresp(split112_merge210_bresp[1:0])
    ,.b_bvalid(split112_merge210_bvalid)
    ,.b_rdata(split112_merge210_rdata[(DWID - 1):0])
    ,.b_rid(split112_merge210_rid[(IDWID - 1):0])
    ,.b_rlast(split112_merge210_rlast)
    ,.b_rready(split112_merge210_rready)
    ,.b_rresp(split112_merge210_rresp[1:0])
    ,.b_rvalid(split112_merge210_rvalid)
    ,.b_wdata(split112_merge210_wdata[(DWID - 1):0])
    ,.b_wlast(split112_merge210_wlast)
    ,.b_wready(split112_merge210_wready)
    ,.b_wstrb(split112_merge210_wstrb[(WSTRB - 1):0])
    ,.b_wvalid(split112_merge210_wvalid)

    ,.c_araddr(split114_merge210_araddr[31:0])
    ,.c_arburst(split114_merge210_arburst[1:0])
    ,.c_arextras(split114_merge210_arextras[(EXTRAS - 1):0])
    ,.c_arid(split114_merge210_arid[(IDWID - 1):0])
    ,.c_arlen(split114_merge210_arlen[7:0])
    ,.c_arready(split114_merge210_arready)
    ,.c_arvalid(split114_merge210_arvalid)
    ,.c_awaddr(split114_merge210_awaddr[31:0])
    ,.c_awburst(split114_merge210_awburst[1:0])
    ,.c_awextras(split114_merge210_awextras[(EXTRAS - 1):0])
    ,.c_awid(split114_merge210_awid[(IDWID - 1):0])
    ,.c_awlen(split114_merge210_awlen[7:0])
    ,.c_awready(split114_merge210_awready)
    ,.c_awvalid(split114_merge210_awvalid)
    ,.c_bid(split114_merge210_bid[(IDWID - 1):0])
    ,.c_bready(split114_merge210_bready)
    ,.c_bresp(split114_merge210_bresp[1:0])
    ,.c_bvalid(split114_merge210_bvalid)
    ,.c_rdata(split114_merge210_rdata[(DWID - 1):0])
    ,.c_rid(split114_merge210_rid[(IDWID - 1):0])
    ,.c_rlast(split114_merge210_rlast)
    ,.c_rready(split114_merge210_rready)
    ,.c_rresp(split114_merge210_rresp[1:0])
    ,.c_rvalid(split114_merge210_rvalid)
    ,.c_wdata(split114_merge210_wdata[(DWID - 1):0])
    ,.c_wlast(split114_merge210_wlast)
    ,.c_wready(split114_merge210_wready)
    ,.c_wstrb(split114_merge210_wstrb[(WSTRB - 1):0])
    ,.c_wvalid(split114_merge210_wvalid)

    ,.d_araddr(split115_merge210_araddr[31:0])
    ,.d_arburst(split115_merge210_arburst[1:0])
    ,.d_arextras(split115_merge210_arextras[(EXTRAS - 1):0])
    ,.d_arid(split115_merge210_arid[(IDWID - 1):0])
    ,.d_arlen(split115_merge210_arlen[7:0])
    ,.d_arready(split115_merge210_arready)
    ,.d_arvalid(split115_merge210_arvalid)
    ,.d_awaddr(split115_merge210_awaddr[31:0])
    ,.d_awburst(split115_merge210_awburst[1:0])
    ,.d_awextras(split115_merge210_awextras[(EXTRAS - 1):0])
    ,.d_awid(split115_merge210_awid[(IDWID - 1):0])
    ,.d_awlen(split115_merge210_awlen[7:0])
    ,.d_awready(split115_merge210_awready)
    ,.d_awvalid(split115_merge210_awvalid)
    ,.d_bid(split115_merge210_bid[(IDWID - 1):0])
    ,.d_bready(split115_merge210_bready)
    ,.d_bresp(split115_merge210_bresp[1:0])
    ,.d_bvalid(split115_merge210_bvalid)
    ,.d_rdata(split115_merge210_rdata[(DWID - 1):0])
    ,.d_rid(split115_merge210_rid[(IDWID - 1):0])
    ,.d_rlast(split115_merge210_rlast)
    ,.d_rready(split115_merge210_rready)
    ,.d_rresp(split115_merge210_rresp[1:0])
    ,.d_rvalid(split115_merge210_rvalid)
    ,.d_wdata(split115_merge210_wdata[(DWID - 1):0])
    ,.d_wlast(split115_merge210_wlast)
    ,.d_wready(split115_merge210_wready)
    ,.d_wstrb(split115_merge210_wstrb[(WSTRB - 1):0])
    ,.d_wvalid(split115_merge210_wvalid)
);


axi_4_merger merge202 (
     .clk(clk),.rst_n(rst_n)
    ,.araddr(slv2_araddr[31:0])
    ,.arburst(slv2_arburst[1:0])
    ,.arextras(slv2_arextras[(EXTRAS - 1):0])
    ,.arid(slv2_arid[(IDWID - 1):0])
    ,.arlen(slv2_arlen[7:0])
    ,.arready(slv2_arready)
    ,.arvalid(slv2_arvalid)
    ,.awaddr(slv2_awaddr[31:0])
    ,.awburst(slv2_awburst[1:0])
    ,.awextras(slv2_awextras[(EXTRAS - 1):0])
    ,.awid(slv2_awid[3:0])
    ,.awlen(slv2_awlen[7:0])
    ,.awready(slv2_awready)
    ,.awvalid(slv2_awvalid)
    ,.bid(slv2_bid[(IDWID - 1):0])
    ,.bready(slv2_bready)
    ,.bresp(slv2_bresp[1:0])
    ,.bvalid(slv2_bvalid)
    ,.rid(slv2_rid[(IDWID - 1):0])
    ,.rlast(slv2_rlast)
    ,.rready(slv2_rready)
    ,.rresp(slv2_rresp[1:0])
    ,.rvalid(slv2_rvalid)
    ,.rdata(slv2_rdata[(DWID - 1):0])
    ,.wdata(slv2_wdata[(DWID - 1):0])
    ,.wlast(slv2_wlast)
    ,.wready(slv2_wready)
    ,.wstrb(slv2_wstrb[(WSTRB - 1):0])
    ,.wvalid(slv2_wvalid)


    ,.a_araddr(split107_merge202_araddr[31:0])
    ,.a_arburst(split107_merge202_arburst[1:0])
    ,.a_arextras(split107_merge202_arextras[(EXTRAS - 1):0])
    ,.a_arid(split107_merge202_arid[(IDWID - 1):0])
    ,.a_arlen(split107_merge202_arlen[7:0])
    ,.a_arready(split107_merge202_arready)
    ,.a_arvalid(split107_merge202_arvalid)
    ,.a_awaddr(split107_merge202_awaddr[31:0])
    ,.a_awburst(split107_merge202_awburst[1:0])
    ,.a_awextras(split107_merge202_awextras[(EXTRAS - 1):0])
    ,.a_awid(split107_merge202_awid[(IDWID - 1):0])
    ,.a_awlen(split107_merge202_awlen[7:0])
    ,.a_awready(split107_merge202_awready)
    ,.a_awvalid(split107_merge202_awvalid)
    ,.a_bid(split107_merge202_bid[(IDWID - 1):0])
    ,.a_bready(split107_merge202_bready)
    ,.a_bresp(split107_merge202_bresp[1:0])
    ,.a_bvalid(split107_merge202_bvalid)
    ,.a_rdata(split107_merge202_rdata[(DWID - 1):0])
    ,.a_rid(split107_merge202_rid[(IDWID - 1):0])
    ,.a_rlast(split107_merge202_rlast)
    ,.a_rready(split107_merge202_rready)
    ,.a_rresp(split107_merge202_rresp[1:0])
    ,.a_rvalid(split107_merge202_rvalid)
    ,.a_wdata(split107_merge202_wdata[(DWID - 1):0])
    ,.a_wlast(split107_merge202_wlast)
    ,.a_wready(split107_merge202_wready)
    ,.a_wstrb(split107_merge202_wstrb[(WSTRB - 1):0])
    ,.a_wvalid(split107_merge202_wvalid)

    ,.b_araddr(split108_merge202_araddr[31:0])
    ,.b_arburst(split108_merge202_arburst[1:0])
    ,.b_arextras(split108_merge202_arextras[(EXTRAS - 1):0])
    ,.b_arid(split108_merge202_arid[(IDWID - 1):0])
    ,.b_arlen(split108_merge202_arlen[7:0])
    ,.b_arready(split108_merge202_arready)
    ,.b_arvalid(split108_merge202_arvalid)
    ,.b_awaddr(split108_merge202_awaddr[31:0])
    ,.b_awburst(split108_merge202_awburst[1:0])
    ,.b_awextras(split108_merge202_awextras[(EXTRAS - 1):0])
    ,.b_awid(split108_merge202_awid[(IDWID - 1):0])
    ,.b_awlen(split108_merge202_awlen[7:0])
    ,.b_awready(split108_merge202_awready)
    ,.b_awvalid(split108_merge202_awvalid)
    ,.b_bid(split108_merge202_bid[(IDWID - 1):0])
    ,.b_bready(split108_merge202_bready)
    ,.b_bresp(split108_merge202_bresp[1:0])
    ,.b_bvalid(split108_merge202_bvalid)
    ,.b_rdata(split108_merge202_rdata[(DWID - 1):0])
    ,.b_rid(split108_merge202_rid[(IDWID - 1):0])
    ,.b_rlast(split108_merge202_rlast)
    ,.b_rready(split108_merge202_rready)
    ,.b_rresp(split108_merge202_rresp[1:0])
    ,.b_rvalid(split108_merge202_rvalid)
    ,.b_wdata(split108_merge202_wdata[(DWID - 1):0])
    ,.b_wlast(split108_merge202_wlast)
    ,.b_wready(split108_merge202_wready)
    ,.b_wstrb(split108_merge202_wstrb[(WSTRB - 1):0])
    ,.b_wvalid(split108_merge202_wvalid)

    ,.c_araddr(split111_merge202_araddr[31:0])
    ,.c_arburst(split111_merge202_arburst[1:0])
    ,.c_arextras(split111_merge202_arextras[(EXTRAS - 1):0])
    ,.c_arid(split111_merge202_arid[(IDWID - 1):0])
    ,.c_arlen(split111_merge202_arlen[7:0])
    ,.c_arready(split111_merge202_arready)
    ,.c_arvalid(split111_merge202_arvalid)
    ,.c_awaddr(split111_merge202_awaddr[31:0])
    ,.c_awburst(split111_merge202_awburst[1:0])
    ,.c_awextras(split111_merge202_awextras[(EXTRAS - 1):0])
    ,.c_awid(split111_merge202_awid[(IDWID - 1):0])
    ,.c_awlen(split111_merge202_awlen[7:0])
    ,.c_awready(split111_merge202_awready)
    ,.c_awvalid(split111_merge202_awvalid)
    ,.c_bid(split111_merge202_bid[(IDWID - 1):0])
    ,.c_bready(split111_merge202_bready)
    ,.c_bresp(split111_merge202_bresp[1:0])
    ,.c_bvalid(split111_merge202_bvalid)
    ,.c_rdata(split111_merge202_rdata[(DWID - 1):0])
    ,.c_rid(split111_merge202_rid[(IDWID - 1):0])
    ,.c_rlast(split111_merge202_rlast)
    ,.c_rready(split111_merge202_rready)
    ,.c_rresp(split111_merge202_rresp[1:0])
    ,.c_rvalid(split111_merge202_rvalid)
    ,.c_wdata(split111_merge202_wdata[(DWID - 1):0])
    ,.c_wlast(split111_merge202_wlast)
    ,.c_wready(split111_merge202_wready)
    ,.c_wstrb(split111_merge202_wstrb[(WSTRB - 1):0])
    ,.c_wvalid(split111_merge202_wvalid)

    ,.d_araddr(split112_merge202_araddr[31:0])
    ,.d_arburst(split112_merge202_arburst[1:0])
    ,.d_arextras(split112_merge202_arextras[(EXTRAS - 1):0])
    ,.d_arid(split112_merge202_arid[(IDWID - 1):0])
    ,.d_arlen(split112_merge202_arlen[7:0])
    ,.d_arready(split112_merge202_arready)
    ,.d_arvalid(split112_merge202_arvalid)
    ,.d_awaddr(split112_merge202_awaddr[31:0])
    ,.d_awburst(split112_merge202_awburst[1:0])
    ,.d_awextras(split112_merge202_awextras[(EXTRAS - 1):0])
    ,.d_awid(split112_merge202_awid[(IDWID - 1):0])
    ,.d_awlen(split112_merge202_awlen[7:0])
    ,.d_awready(split112_merge202_awready)
    ,.d_awvalid(split112_merge202_awvalid)
    ,.d_bid(split112_merge202_bid[(IDWID - 1):0])
    ,.d_bready(split112_merge202_bready)
    ,.d_bresp(split112_merge202_bresp[1:0])
    ,.d_bvalid(split112_merge202_bvalid)
    ,.d_rdata(split112_merge202_rdata[(DWID - 1):0])
    ,.d_rid(split112_merge202_rid[(IDWID - 1):0])
    ,.d_rlast(split112_merge202_rlast)
    ,.d_rready(split112_merge202_rready)
    ,.d_rresp(split112_merge202_rresp[1:0])
    ,.d_rvalid(split112_merge202_rvalid)
    ,.d_wdata(split112_merge202_wdata[(DWID - 1):0])
    ,.d_wlast(split112_merge202_wlast)
    ,.d_wready(split112_merge202_wready)
    ,.d_wstrb(split112_merge202_wstrb[(WSTRB - 1):0])
    ,.d_wvalid(split112_merge202_wvalid)
);


axi_4_merger merge215 (
     .clk(clk),.rst_n(rst_n)
    ,.araddr(slv15_araddr[31:0])
    ,.arburst(slv15_arburst[1:0])
    ,.arextras(slv15_arextras[(EXTRAS - 1):0])
    ,.arid(slv15_arid[(IDWID - 1):0])
    ,.arlen(slv15_arlen[7:0])
    ,.arready(slv15_arready)
    ,.arvalid(slv15_arvalid)
    ,.awaddr(slv15_awaddr[31:0])
    ,.awburst(slv15_awburst[1:0])
    ,.awextras(slv15_awextras[(EXTRAS - 1):0])
    ,.awid(slv15_awid[3:0])
    ,.awlen(slv15_awlen[7:0])
    ,.awready(slv15_awready)
    ,.awvalid(slv15_awvalid)
    ,.bid(slv15_bid[(IDWID - 1):0])
    ,.bready(slv15_bready)
    ,.bresp(slv15_bresp[1:0])
    ,.bvalid(slv15_bvalid)
    ,.rid(slv15_rid[(IDWID - 1):0])
    ,.rlast(slv15_rlast)
    ,.rready(slv15_rready)
    ,.rresp(slv15_rresp[1:0])
    ,.rvalid(slv15_rvalid)
    ,.rdata(slv15_rdata[(DWID - 1):0])
    ,.wdata(slv15_wdata[(DWID - 1):0])
    ,.wlast(slv15_wlast)
    ,.wready(slv15_wready)
    ,.wstrb(slv15_wstrb[(WSTRB - 1):0])
    ,.wvalid(slv15_wvalid)


    ,.a_araddr(split109_merge215_araddr[31:0])
    ,.a_arburst(split109_merge215_arburst[1:0])
    ,.a_arextras(split109_merge215_arextras[(EXTRAS - 1):0])
    ,.a_arid(split109_merge215_arid[(IDWID - 1):0])
    ,.a_arlen(split109_merge215_arlen[7:0])
    ,.a_arready(split109_merge215_arready)
    ,.a_arvalid(split109_merge215_arvalid)
    ,.a_awaddr(split109_merge215_awaddr[31:0])
    ,.a_awburst(split109_merge215_awburst[1:0])
    ,.a_awextras(split109_merge215_awextras[(EXTRAS - 1):0])
    ,.a_awid(split109_merge215_awid[(IDWID - 1):0])
    ,.a_awlen(split109_merge215_awlen[7:0])
    ,.a_awready(split109_merge215_awready)
    ,.a_awvalid(split109_merge215_awvalid)
    ,.a_bid(split109_merge215_bid[(IDWID - 1):0])
    ,.a_bready(split109_merge215_bready)
    ,.a_bresp(split109_merge215_bresp[1:0])
    ,.a_bvalid(split109_merge215_bvalid)
    ,.a_rdata(split109_merge215_rdata[(DWID - 1):0])
    ,.a_rid(split109_merge215_rid[(IDWID - 1):0])
    ,.a_rlast(split109_merge215_rlast)
    ,.a_rready(split109_merge215_rready)
    ,.a_rresp(split109_merge215_rresp[1:0])
    ,.a_rvalid(split109_merge215_rvalid)
    ,.a_wdata(split109_merge215_wdata[(DWID - 1):0])
    ,.a_wlast(split109_merge215_wlast)
    ,.a_wready(split109_merge215_wready)
    ,.a_wstrb(split109_merge215_wstrb[(WSTRB - 1):0])
    ,.a_wvalid(split109_merge215_wvalid)

    ,.b_araddr(split110_merge215_araddr[31:0])
    ,.b_arburst(split110_merge215_arburst[1:0])
    ,.b_arextras(split110_merge215_arextras[(EXTRAS - 1):0])
    ,.b_arid(split110_merge215_arid[(IDWID - 1):0])
    ,.b_arlen(split110_merge215_arlen[7:0])
    ,.b_arready(split110_merge215_arready)
    ,.b_arvalid(split110_merge215_arvalid)
    ,.b_awaddr(split110_merge215_awaddr[31:0])
    ,.b_awburst(split110_merge215_awburst[1:0])
    ,.b_awextras(split110_merge215_awextras[(EXTRAS - 1):0])
    ,.b_awid(split110_merge215_awid[(IDWID - 1):0])
    ,.b_awlen(split110_merge215_awlen[7:0])
    ,.b_awready(split110_merge215_awready)
    ,.b_awvalid(split110_merge215_awvalid)
    ,.b_bid(split110_merge215_bid[(IDWID - 1):0])
    ,.b_bready(split110_merge215_bready)
    ,.b_bresp(split110_merge215_bresp[1:0])
    ,.b_bvalid(split110_merge215_bvalid)
    ,.b_rdata(split110_merge215_rdata[(DWID - 1):0])
    ,.b_rid(split110_merge215_rid[(IDWID - 1):0])
    ,.b_rlast(split110_merge215_rlast)
    ,.b_rready(split110_merge215_rready)
    ,.b_rresp(split110_merge215_rresp[1:0])
    ,.b_rvalid(split110_merge215_rvalid)
    ,.b_wdata(split110_merge215_wdata[(DWID - 1):0])
    ,.b_wlast(split110_merge215_wlast)
    ,.b_wready(split110_merge215_wready)
    ,.b_wstrb(split110_merge215_wstrb[(WSTRB - 1):0])
    ,.b_wvalid(split110_merge215_wvalid)

    ,.c_araddr(split112_merge215_araddr[31:0])
    ,.c_arburst(split112_merge215_arburst[1:0])
    ,.c_arextras(split112_merge215_arextras[(EXTRAS - 1):0])
    ,.c_arid(split112_merge215_arid[(IDWID - 1):0])
    ,.c_arlen(split112_merge215_arlen[7:0])
    ,.c_arready(split112_merge215_arready)
    ,.c_arvalid(split112_merge215_arvalid)
    ,.c_awaddr(split112_merge215_awaddr[31:0])
    ,.c_awburst(split112_merge215_awburst[1:0])
    ,.c_awextras(split112_merge215_awextras[(EXTRAS - 1):0])
    ,.c_awid(split112_merge215_awid[(IDWID - 1):0])
    ,.c_awlen(split112_merge215_awlen[7:0])
    ,.c_awready(split112_merge215_awready)
    ,.c_awvalid(split112_merge215_awvalid)
    ,.c_bid(split112_merge215_bid[(IDWID - 1):0])
    ,.c_bready(split112_merge215_bready)
    ,.c_bresp(split112_merge215_bresp[1:0])
    ,.c_bvalid(split112_merge215_bvalid)
    ,.c_rdata(split112_merge215_rdata[(DWID - 1):0])
    ,.c_rid(split112_merge215_rid[(IDWID - 1):0])
    ,.c_rlast(split112_merge215_rlast)
    ,.c_rready(split112_merge215_rready)
    ,.c_rresp(split112_merge215_rresp[1:0])
    ,.c_rvalid(split112_merge215_rvalid)
    ,.c_wdata(split112_merge215_wdata[(DWID - 1):0])
    ,.c_wlast(split112_merge215_wlast)
    ,.c_wready(split112_merge215_wready)
    ,.c_wstrb(split112_merge215_wstrb[(WSTRB - 1):0])
    ,.c_wvalid(split112_merge215_wvalid)

    ,.d_araddr(split114_merge215_araddr[31:0])
    ,.d_arburst(split114_merge215_arburst[1:0])
    ,.d_arextras(split114_merge215_arextras[(EXTRAS - 1):0])
    ,.d_arid(split114_merge215_arid[(IDWID - 1):0])
    ,.d_arlen(split114_merge215_arlen[7:0])
    ,.d_arready(split114_merge215_arready)
    ,.d_arvalid(split114_merge215_arvalid)
    ,.d_awaddr(split114_merge215_awaddr[31:0])
    ,.d_awburst(split114_merge215_awburst[1:0])
    ,.d_awextras(split114_merge215_awextras[(EXTRAS - 1):0])
    ,.d_awid(split114_merge215_awid[(IDWID - 1):0])
    ,.d_awlen(split114_merge215_awlen[7:0])
    ,.d_awready(split114_merge215_awready)
    ,.d_awvalid(split114_merge215_awvalid)
    ,.d_bid(split114_merge215_bid[(IDWID - 1):0])
    ,.d_bready(split114_merge215_bready)
    ,.d_bresp(split114_merge215_bresp[1:0])
    ,.d_bvalid(split114_merge215_bvalid)
    ,.d_rdata(split114_merge215_rdata[(DWID - 1):0])
    ,.d_rid(split114_merge215_rid[(IDWID - 1):0])
    ,.d_rlast(split114_merge215_rlast)
    ,.d_rready(split114_merge215_rready)
    ,.d_rresp(split114_merge215_rresp[1:0])
    ,.d_rvalid(split114_merge215_rvalid)
    ,.d_wdata(split114_merge215_wdata[(DWID - 1):0])
    ,.d_wlast(split114_merge215_wlast)
    ,.d_wready(split114_merge215_wready)
    ,.d_wstrb(split114_merge215_wstrb[(WSTRB - 1):0])
    ,.d_wvalid(split114_merge215_wvalid)
);



reg [1023:0] testname;
initial begin
   if ($value$plusargs("LOG=%s",testname)) begin 
        $python("pymonname()",testname);
    end  


    if ($value$plusargs("SEQ=%s",testname)) begin 
         $display(" Running SEQ= %s.",testname); 
    end else begin
        testname = 0; 
        $display(" default test");
    end  
    #10; 
    if (testname!=0) $python("sequence()",testname);
end 
endmodule

