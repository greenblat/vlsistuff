`define DEMO_BASEADDR    'h0
`define ADDR_KEY0                                                'h0
`define ADDR_KEY1                                                'h10
`define ADDR_LIMITS0                                             'h20
`define ADDR_LIMITS1                                             'h40
