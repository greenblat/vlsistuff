module smalltab (input [9:0] ain, output [31:0] out);
assign out = 
    (ain==1) ? 32'h3f801630 :
    (ain==2) ? 32'h3f802c64 :
    (ain==3) ? 32'h3f80429c :
    (ain==4) ? 32'h3f8058d7 :
    (ain==5) ? 32'h3f806f17 :
    (ain==6) ? 32'h3f80855a :
    (ain==7) ? 32'h3f809ba2 :
    (ain==8) ? 32'h3f80b1ed :
    (ain==9) ? 32'h3f80c83c :
    (ain==10) ? 32'h3f80de8f :
    (ain==11) ? 32'h3f80f4e5 :
    (ain==12) ? 32'h3f810b40 :
    (ain==13) ? 32'h3f81219f :
    (ain==14) ? 32'h3f813801 :
    (ain==15) ? 32'h3f814e67 :
    (ain==16) ? 32'h3f8164d1 :
    (ain==17) ? 32'h3f817b3f :
    (ain==18) ? 32'h3f8191b1 :
    (ain==19) ? 32'h3f81a827 :
    (ain==20) ? 32'h3f81bea1 :
    (ain==21) ? 32'h3f81d51f :
    (ain==22) ? 32'h3f81eba0 :
    (ain==23) ? 32'h3f820225 :
    (ain==24) ? 32'h3f8218af :
    (ain==25) ? 32'h3f822f3c :
    (ain==26) ? 32'h3f8245cd :
    (ain==27) ? 32'h3f825c62 :
    (ain==28) ? 32'h3f8272fb :
    (ain==29) ? 32'h3f828998 :
    (ain==30) ? 32'h3f82a039 :
    (ain==31) ? 32'h3f82b6dd :
    (ain==32) ? 32'h3f82cd86 :
    (ain==33) ? 32'h3f82e433 :
    (ain==34) ? 32'h3f82fae3 :
    (ain==35) ? 32'h3f831198 :
    (ain==36) ? 32'h3f832850 :
    (ain==37) ? 32'h3f833f0c :
    (ain==38) ? 32'h3f8355cc :
    (ain==39) ? 32'h3f836c91 :
    (ain==40) ? 32'h3f838359 :
    (ain==41) ? 32'h3f839a25 :
    (ain==42) ? 32'h3f83b0f5 :
    (ain==43) ? 32'h3f83c7c9 :
    (ain==44) ? 32'h3f83dea1 :
    (ain==45) ? 32'h3f83f57d :
    (ain==46) ? 32'h3f840c5d :
    (ain==47) ? 32'h3f842340 :
    (ain==48) ? 32'h3f843a28 :
    (ain==49) ? 32'h3f845114 :
    (ain==50) ? 32'h3f846804 :
    (ain==51) ? 32'h3f847ef8 :
    (ain==52) ? 32'h3f8495ef :
    (ain==53) ? 32'h3f84aceb :
    (ain==54) ? 32'h3f84c3eb :
    (ain==55) ? 32'h3f84daee :
    (ain==56) ? 32'h3f84f1f6 :
    (ain==57) ? 32'h3f850901 :
    (ain==58) ? 32'h3f852011 :
    (ain==59) ? 32'h3f853725 :
    (ain==60) ? 32'h3f854e3c :
    (ain==61) ? 32'h3f856558 :
    (ain==62) ? 32'h3f857c78 :
    (ain==63) ? 32'h3f85939b :
    (ain==64) ? 32'h3f85aac3 :
    (ain==65) ? 32'h3f85c1ef :
    (ain==66) ? 32'h3f85d91e :
    (ain==67) ? 32'h3f85f052 :
    (ain==68) ? 32'h3f86078a :
    (ain==69) ? 32'h3f861ec5 :
    (ain==70) ? 32'h3f863605 :
    (ain==71) ? 32'h3f864d49 :
    (ain==72) ? 32'h3f866491 :
    (ain==73) ? 32'h3f867bdd :
    (ain==74) ? 32'h3f86932d :
    (ain==75) ? 32'h3f86aa81 :
    (ain==76) ? 32'h3f86c1d9 :
    (ain==77) ? 32'h3f86d935 :
    (ain==78) ? 32'h3f86f095 :
    (ain==79) ? 32'h3f8707f9 :
    (ain==80) ? 32'h3f871f61 :
    (ain==81) ? 32'h3f8736cd :
    (ain==82) ? 32'h3f874e3e :
    (ain==83) ? 32'h3f8765b2 :
    (ain==84) ? 32'h3f877d2a :
    (ain==85) ? 32'h3f8794a7 :
    (ain==86) ? 32'h3f87ac28 :
    (ain==87) ? 32'h3f87c3ac :
    (ain==88) ? 32'h3f87db35 :
    (ain==89) ? 32'h3f87f2c2 :
    (ain==90) ? 32'h3f880a53 :
    (ain==91) ? 32'h3f8821e8 :
    (ain==92) ? 32'h3f883981 :
    (ain==93) ? 32'h3f88511e :
    (ain==94) ? 32'h3f8868bf :
    (ain==95) ? 32'h3f888065 :
    (ain==96) ? 32'h3f88980e :
    (ain==97) ? 32'h3f88afbc :
    (ain==98) ? 32'h3f88c76d :
    (ain==99) ? 32'h3f88df23 :
    (ain==100) ? 32'h3f88f6dd :
    (ain==101) ? 32'h3f890e9b :
    (ain==102) ? 32'h3f89265d :
    (ain==103) ? 32'h3f893e23 :
    (ain==104) ? 32'h3f8955ee :
    (ain==105) ? 32'h3f896dbc :
    (ain==106) ? 32'h3f89858f :
    (ain==107) ? 32'h3f899d65 :
    (ain==108) ? 32'h3f89b540 :
    (ain==109) ? 32'h3f89cd1f :
    (ain==110) ? 32'h3f89e502 :
    (ain==111) ? 32'h3f89fcea :
    (ain==112) ? 32'h3f8a14d5 :
    (ain==113) ? 32'h3f8a2cc5 :
    (ain==114) ? 32'h3f8a44b8 :
    (ain==115) ? 32'h3f8a5cb0 :
    (ain==116) ? 32'h3f8a74ac :
    (ain==117) ? 32'h3f8a8cac :
    (ain==118) ? 32'h3f8aa4b1 :
    (ain==119) ? 32'h3f8abcb9 :
    (ain==120) ? 32'h3f8ad4c6 :
    (ain==121) ? 32'h3f8aecd7 :
    (ain==122) ? 32'h3f8b04ec :
    (ain==123) ? 32'h3f8b1d05 :
    (ain==124) ? 32'h3f8b3522 :
    (ain==125) ? 32'h3f8b4d44 :
    (ain==126) ? 32'h3f8b6569 :
    (ain==127) ? 32'h3f8b7d93 :
    (ain==128) ? 32'h3f8b95c1 :
    (ain==129) ? 32'h3f8badf4 :
    (ain==130) ? 32'h3f8bc62a :
    (ain==131) ? 32'h3f8bde65 :
    (ain==132) ? 32'h3f8bf6a4 :
    (ain==133) ? 32'h3f8c0ee7 :
    (ain==134) ? 32'h3f8c272e :
    (ain==135) ? 32'h3f8c3f7a :
    (ain==136) ? 32'h3f8c57c9 :
    (ain==137) ? 32'h3f8c701d :
    (ain==138) ? 32'h3f8c8875 :
    (ain==139) ? 32'h3f8ca0d2 :
    (ain==140) ? 32'h3f8cb932 :
    (ain==141) ? 32'h3f8cd197 :
    (ain==142) ? 32'h3f8cea00 :
    (ain==143) ? 32'h3f8d026d :
    (ain==144) ? 32'h3f8d1adf :
    (ain==145) ? 32'h3f8d3355 :
    (ain==146) ? 32'h3f8d4bcf :
    (ain==147) ? 32'h3f8d644d :
    (ain==148) ? 32'h3f8d7ccf :
    (ain==149) ? 32'h3f8d9556 :
    (ain==150) ? 32'h3f8dade1 :
    (ain==151) ? 32'h3f8dc670 :
    (ain==152) ? 32'h3f8ddf04 :
    (ain==153) ? 32'h3f8df79b :
    (ain==154) ? 32'h3f8e1037 :
    (ain==155) ? 32'h3f8e28d8 :
    (ain==156) ? 32'h3f8e417c :
    (ain==157) ? 32'h3f8e5a25 :
    (ain==158) ? 32'h3f8e72d2 :
    (ain==159) ? 32'h3f8e8b83 :
    (ain==160) ? 32'h3f8ea439 :
    (ain==161) ? 32'h3f8ebcf3 :
    (ain==162) ? 32'h3f8ed5b1 :
    (ain==163) ? 32'h3f8eee74 :
    (ain==164) ? 32'h3f8f073a :
    (ain==165) ? 32'h3f8f2006 :
    (ain==166) ? 32'h3f8f38d5 :
    (ain==167) ? 32'h3f8f51a9 :
    (ain==168) ? 32'h3f8f6a81 :
    (ain==169) ? 32'h3f8f835d :
    (ain==170) ? 32'h3f8f9c3d :
    (ain==171) ? 32'h3f8fb522 :
    (ain==172) ? 32'h3f8fce0c :
    (ain==173) ? 32'h3f8fe6f9 :
    (ain==174) ? 32'h3f8fffeb :
    (ain==175) ? 32'h3f9018e1 :
    (ain==176) ? 32'h3f9031dc :
    (ain==177) ? 32'h3f904adb :
    (ain==178) ? 32'h3f9063de :
    (ain==179) ? 32'h3f907ce5 :
    (ain==180) ? 32'h3f9095f1 :
    (ain==181) ? 32'h3f90af01 :
    (ain==182) ? 32'h3f90c816 :
    (ain==183) ? 32'h3f90e12f :
    (ain==184) ? 32'h3f90fa4c :
    (ain==185) ? 32'h3f91136e :
    (ain==186) ? 32'h3f912c94 :
    (ain==187) ? 32'h3f9145be :
    (ain==188) ? 32'h3f915eed :
    (ain==189) ? 32'h3f917820 :
    (ain==190) ? 32'h3f919157 :
    (ain==191) ? 32'h3f91aa93 :
    (ain==192) ? 32'h3f91c3d3 :
    (ain==193) ? 32'h3f91dd17 :
    (ain==194) ? 32'h3f91f660 :
    (ain==195) ? 32'h3f920fae :
    (ain==196) ? 32'h3f9228ff :
    (ain==197) ? 32'h3f924255 :
    (ain==198) ? 32'h3f925bb0 :
    (ain==199) ? 32'h3f92750f :
    (ain==200) ? 32'h3f928e72 :
    (ain==201) ? 32'h3f92a7da :
    (ain==202) ? 32'h3f92c146 :
    (ain==203) ? 32'h3f92dab6 :
    (ain==204) ? 32'h3f92f42b :
    (ain==205) ? 32'h3f930da4 :
    (ain==206) ? 32'h3f932722 :
    (ain==207) ? 32'h3f9340a4 :
    (ain==208) ? 32'h3f935a2b :
    (ain==209) ? 32'h3f9373b6 :
    (ain==210) ? 32'h3f938d45 :
    (ain==211) ? 32'h3f93a6d9 :
    (ain==212) ? 32'h3f93c071 :
    (ain==213) ? 32'h3f93da0e :
    (ain==214) ? 32'h3f93f3af :
    (ain==215) ? 32'h3f940d55 :
    (ain==216) ? 32'h3f9426ff :
    (ain==217) ? 32'h3f9440ad :
    (ain==218) ? 32'h3f945a60 :
    (ain==219) ? 32'h3f947417 :
    (ain==220) ? 32'h3f948dd3 :
    (ain==221) ? 32'h3f94a793 :
    (ain==222) ? 32'h3f94c158 :
    (ain==223) ? 32'h3f94db21 :
    (ain==224) ? 32'h3f94f4ef :
    (ain==225) ? 32'h3f950ec1 :
    (ain==226) ? 32'h3f952898 :
    (ain==227) ? 32'h3f954273 :
    (ain==228) ? 32'h3f955c53 :
    (ain==229) ? 32'h3f957637 :
    (ain==230) ? 32'h3f95901f :
    (ain==231) ? 32'h3f95aa0c :
    (ain==232) ? 32'h3f95c3fe :
    (ain==233) ? 32'h3f95ddf4 :
    (ain==234) ? 32'h3f95f7ef :
    (ain==235) ? 32'h3f9611ee :
    (ain==236) ? 32'h3f962bf1 :
    (ain==237) ? 32'h3f9645f9 :
    (ain==238) ? 32'h3f966006 :
    (ain==239) ? 32'h3f967a17 :
    (ain==240) ? 32'h3f96942d :
    (ain==241) ? 32'h3f96ae47 :
    (ain==242) ? 32'h3f96c866 :
    (ain==243) ? 32'h3f96e289 :
    (ain==244) ? 32'h3f96fcb0 :
    (ain==245) ? 32'h3f9716dd :
    (ain==246) ? 32'h3f97310e :
    (ain==247) ? 32'h3f974b43 :
    (ain==248) ? 32'h3f97657d :
    (ain==249) ? 32'h3f977fbb :
    (ain==250) ? 32'h3f9799fe :
    (ain==251) ? 32'h3f97b446 :
    (ain==252) ? 32'h3f97ce92 :
    (ain==253) ? 32'h3f97e8e2 :
    (ain==254) ? 32'h3f980338 :
    (ain==255) ? 32'h3f981d91 :
    (ain==256) ? 32'h3f9837f0 :
    (ain==257) ? 32'h3f985253 :
    (ain==258) ? 32'h3f986cba :
    (ain==259) ? 32'h3f988726 :
    (ain==260) ? 32'h3f98a197 :
    (ain==261) ? 32'h3f98bc0c :
    (ain==262) ? 32'h3f98d686 :
    (ain==263) ? 32'h3f98f104 :
    (ain==264) ? 32'h3f990b87 :
    (ain==265) ? 32'h3f99260f :
    (ain==266) ? 32'h3f99409b :
    (ain==267) ? 32'h3f995b2c :
    (ain==268) ? 32'h3f9975c1 :
    (ain==269) ? 32'h3f99905b :
    (ain==270) ? 32'h3f99aafa :
    (ain==271) ? 32'h3f99c59d :
    (ain==272) ? 32'h3f99e045 :
    (ain==273) ? 32'h3f99faf2 :
    (ain==274) ? 32'h3f9a15a3 :
    (ain==275) ? 32'h3f9a3058 :
    (ain==276) ? 32'h3f9a4b13 :
    (ain==277) ? 32'h3f9a65d2 :
    (ain==278) ? 32'h3f9a8095 :
    (ain==279) ? 32'h3f9a9b5e :
    (ain==280) ? 32'h3f9ab62a :
    (ain==281) ? 32'h3f9ad0fc :
    (ain==282) ? 32'h3f9aebd2 :
    (ain==283) ? 32'h3f9b06ad :
    (ain==284) ? 32'h3f9b218d :
    (ain==285) ? 32'h3f9b3c71 :
    (ain==286) ? 32'h3f9b575a :
    (ain==287) ? 32'h3f9b7247 :
    (ain==288) ? 32'h3f9b8d39 :
    (ain==289) ? 32'h3f9ba830 :
    (ain==290) ? 32'h3f9bc32c :
    (ain==291) ? 32'h3f9bde2c :
    (ain==292) ? 32'h3f9bf931 :
    (ain==293) ? 32'h3f9c143a :
    (ain==294) ? 32'h3f9c2f48 :
    (ain==295) ? 32'h3f9c4a5b :
    (ain==296) ? 32'h3f9c6573 :
    (ain==297) ? 32'h3f9c808f :
    (ain==298) ? 32'h3f9c9bb0 :
    (ain==299) ? 32'h3f9cb6d6 :
    (ain==300) ? 32'h3f9cd200 :
    (ain==301) ? 32'h3f9ced2f :
    (ain==302) ? 32'h3f9d0863 :
    (ain==303) ? 32'h3f9d239c :
    (ain==304) ? 32'h3f9d3ed9 :
    (ain==305) ? 32'h3f9d5a1b :
    (ain==306) ? 32'h3f9d7562 :
    (ain==307) ? 32'h3f9d90ad :
    (ain==308) ? 32'h3f9dabfd :
    (ain==309) ? 32'h3f9dc752 :
    (ain==310) ? 32'h3f9de2ac :
    (ain==311) ? 32'h3f9dfe0a :
    (ain==312) ? 32'h3f9e196e :
    (ain==313) ? 32'h3f9e34d5 :
    (ain==314) ? 32'h3f9e5042 :
    (ain==315) ? 32'h3f9e6bb4 :
    (ain==316) ? 32'h3f9e872a :
    (ain==317) ? 32'h3f9ea2a5 :
    (ain==318) ? 32'h3f9ebe24 :
    (ain==319) ? 32'h3f9ed9a9 :
    (ain==320) ? 32'h3f9ef532 :
    (ain==321) ? 32'h3f9f10c0 :
    (ain==322) ? 32'h3f9f2c53 :
    (ain==323) ? 32'h3f9f47ea :
    (ain==324) ? 32'h3f9f6386 :
    (ain==325) ? 32'h3f9f7f28 :
    (ain==326) ? 32'h3f9f9acd :
    (ain==327) ? 32'h3f9fb678 :
    (ain==328) ? 32'h3f9fd228 :
    (ain==329) ? 32'h3f9feddc :
    (ain==330) ? 32'h3fa00995 :
    (ain==331) ? 32'h3fa02553 :
    (ain==332) ? 32'h3fa04116 :
    (ain==333) ? 32'h3fa05cdd :
    (ain==334) ? 32'h3fa078a9 :
    (ain==335) ? 32'h3fa0947b :
    (ain==336) ? 32'h3fa0b051 :
    (ain==337) ? 32'h3fa0cc2b :
    (ain==338) ? 32'h3fa0e80b :
    (ain==339) ? 32'h3fa103ef :
    (ain==340) ? 32'h3fa11fd9 :
    (ain==341) ? 32'h3fa13bc7 :
    (ain==342) ? 32'h3fa157ba :
    (ain==343) ? 32'h3fa173b2 :
    (ain==344) ? 32'h3fa18fae :
    (ain==345) ? 32'h3fa1abb0 :
    (ain==346) ? 32'h3fa1c7b6 :
    (ain==347) ? 32'h3fa1e3c1 :
    (ain==348) ? 32'h3fa1ffd1 :
    (ain==349) ? 32'h3fa21be6 :
    (ain==350) ? 32'h3fa23800 :
    (ain==351) ? 32'h3fa2541f :
    (ain==352) ? 32'h3fa27043 :
    (ain==353) ? 32'h3fa28c6b :
    (ain==354) ? 32'h3fa2a898 :
    (ain==355) ? 32'h3fa2c4ca :
    (ain==356) ? 32'h3fa2e102 :
    (ain==357) ? 32'h3fa2fd3e :
    (ain==358) ? 32'h3fa3197e :
    (ain==359) ? 32'h3fa335c4 :
    (ain==360) ? 32'h3fa3520f :
    (ain==361) ? 32'h3fa36e5e :
    (ain==362) ? 32'h3fa38ab3 :
    (ain==363) ? 32'h3fa3a70c :
    (ain==364) ? 32'h3fa3c36b :
    (ain==365) ? 32'h3fa3dfce :
    (ain==366) ? 32'h3fa3fc36 :
    (ain==367) ? 32'h3fa418a3 :
    (ain==368) ? 32'h3fa43515 :
    (ain==369) ? 32'h3fa4518c :
    (ain==370) ? 32'h3fa46e08 :
    (ain==371) ? 32'h3fa48a89 :
    (ain==372) ? 32'h3fa4a70f :
    (ain==373) ? 32'h3fa4c399 :
    (ain==374) ? 32'h3fa4e029 :
    (ain==375) ? 32'h3fa4fcbd :
    (ain==376) ? 32'h3fa51957 :
    (ain==377) ? 32'h3fa535f6 :
    (ain==378) ? 32'h3fa55299 :
    (ain==379) ? 32'h3fa56f41 :
    (ain==380) ? 32'h3fa58bef :
    (ain==381) ? 32'h3fa5a8a1 :
    (ain==382) ? 32'h3fa5c559 :
    (ain==383) ? 32'h3fa5e215 :
    (ain==384) ? 32'h3fa5fed6 :
    (ain==385) ? 32'h3fa61b9c :
    (ain==386) ? 32'h3fa63868 :
    (ain==387) ? 32'h3fa65538 :
    (ain==388) ? 32'h3fa6720d :
    (ain==389) ? 32'h3fa68ee8 :
    (ain==390) ? 32'h3fa6abc7 :
    (ain==391) ? 32'h3fa6c8ab :
    (ain==392) ? 32'h3fa6e594 :
    (ain==393) ? 32'h3fa70283 :
    (ain==394) ? 32'h3fa71f76 :
    (ain==395) ? 32'h3fa73c6e :
    (ain==396) ? 32'h3fa7596c :
    (ain==397) ? 32'h3fa7766e :
    (ain==398) ? 32'h3fa79375 :
    (ain==399) ? 32'h3fa7b082 :
    (ain==400) ? 32'h3fa7cd93 :
    (ain==401) ? 32'h3fa7eaaa :
    (ain==402) ? 32'h3fa807c5 :
    (ain==403) ? 32'h3fa824e6 :
    (ain==404) ? 32'h3fa8420b :
    (ain==405) ? 32'h3fa85f36 :
    (ain==406) ? 32'h3fa87c66 :
    (ain==407) ? 32'h3fa8999b :
    (ain==408) ? 32'h3fa8b6d5 :
    (ain==409) ? 32'h3fa8d414 :
    (ain==410) ? 32'h3fa8f158 :
    (ain==411) ? 32'h3fa90ea1 :
    (ain==412) ? 32'h3fa92bef :
    (ain==413) ? 32'h3fa94942 :
    (ain==414) ? 32'h3fa9669a :
    (ain==415) ? 32'h3fa983f8 :
    (ain==416) ? 32'h3fa9a15a :
    (ain==417) ? 32'h3fa9bec2 :
    (ain==418) ? 32'h3fa9dc2e :
    (ain==419) ? 32'h3fa9f9a0 :
    (ain==420) ? 32'h3faa1717 :
    (ain==421) ? 32'h3faa3493 :
    (ain==422) ? 32'h3faa5214 :
    (ain==423) ? 32'h3faa6f9a :
    (ain==424) ? 32'h3faa8d26 :
    (ain==425) ? 32'h3faaaab6 :
    (ain==426) ? 32'h3faac84c :
    (ain==427) ? 32'h3faae5e7 :
    (ain==428) ? 32'h3fab0386 :
    (ain==429) ? 32'h3fab212b :
    (ain==430) ? 32'h3fab3ed6 :
    (ain==431) ? 32'h3fab5c85 :
    (ain==432) ? 32'h3fab7a39 :
    (ain==433) ? 32'h3fab97f3 :
    (ain==434) ? 32'h3fabb5b1 :
    (ain==435) ? 32'h3fabd375 :
    (ain==436) ? 32'h3fabf13e :
    (ain==437) ? 32'h3fac0f0d :
    (ain==438) ? 32'h3fac2ce0 :
    (ain==439) ? 32'h3fac4ab8 :
    (ain==440) ? 32'h3fac6896 :
    (ain==441) ? 32'h3fac8679 :
    (ain==442) ? 32'h3faca461 :
    (ain==443) ? 32'h3facc24e :
    (ain==444) ? 32'h3face041 :
    (ain==445) ? 32'h3facfe38 :
    (ain==446) ? 32'h3fad1c35 :
    (ain==447) ? 32'h3fad3a37 :
    (ain==448) ? 32'h3fad583e :
    (ain==449) ? 32'h3fad764b :
    (ain==450) ? 32'h3fad945c :
    (ain==451) ? 32'h3fadb273 :
    (ain==452) ? 32'h3fadd08f :
    (ain==453) ? 32'h3fadeeb1 :
    (ain==454) ? 32'h3fae0cd7 :
    (ain==455) ? 32'h3fae2b03 :
    (ain==456) ? 32'h3fae4934 :
    (ain==457) ? 32'h3fae676a :
    (ain==458) ? 32'h3fae85a5 :
    (ain==459) ? 32'h3faea3e6 :
    (ain==460) ? 32'h3faec22c :
    (ain==461) ? 32'h3faee077 :
    (ain==462) ? 32'h3faefec8 :
    (ain==463) ? 32'h3faf1d1d :
    (ain==464) ? 32'h3faf3b78 :
    (ain==465) ? 32'h3faf59d8 :
    (ain==466) ? 32'h3faf783e :
    (ain==467) ? 32'h3faf96a9 :
    (ain==468) ? 32'h3fafb519 :
    (ain==469) ? 32'h3fafd38e :
    (ain==470) ? 32'h3faff208 :
    (ain==471) ? 32'h3fb01088 :
    (ain==472) ? 32'h3fb02f0d :
    (ain==473) ? 32'h3fb04d98 :
    (ain==474) ? 32'h3fb06c27 :
    (ain==475) ? 32'h3fb08abc :
    (ain==476) ? 32'h3fb0a957 :
    (ain==477) ? 32'h3fb0c7f6 :
    (ain==478) ? 32'h3fb0e69b :
    (ain==479) ? 32'h3fb10545 :
    (ain==480) ? 32'h3fb123f5 :
    (ain==481) ? 32'h3fb142aa :
    (ain==482) ? 32'h3fb16164 :
    (ain==483) ? 32'h3fb18024 :
    (ain==484) ? 32'h3fb19ee8 :
    (ain==485) ? 32'h3fb1bdb3 :
    (ain==486) ? 32'h3fb1dc82 :
    (ain==487) ? 32'h3fb1fb57 :
    (ain==488) ? 32'h3fb21a31 :
    (ain==489) ? 32'h3fb23911 :
    (ain==490) ? 32'h3fb257f6 :
    (ain==491) ? 32'h3fb276e0 :
    (ain==492) ? 32'h3fb295cf :
    (ain==493) ? 32'h3fb2b4c4 :
    (ain==494) ? 32'h3fb2d3bf :
    (ain==495) ? 32'h3fb2f2be :
    (ain==496) ? 32'h3fb311c4 :
    (ain==497) ? 32'h3fb330ce :
    (ain==498) ? 32'h3fb34fde :
    (ain==499) ? 32'h3fb36ef3 :
    (ain==500) ? 32'h3fb38e0e :
    (ain==501) ? 32'h3fb3ad2e :
    (ain==502) ? 32'h3fb3cc53 :
    (ain==503) ? 32'h3fb3eb7e :
    (ain==504) ? 32'h3fb40aae :
    (ain==505) ? 32'h3fb429e4 :
    (ain==506) ? 32'h3fb4491f :
    (ain==507) ? 32'h3fb4685f :
    (ain==508) ? 32'h3fb487a5 :
    (ain==509) ? 32'h3fb4a6f0 :
    (ain==510) ? 32'h3fb4c641 :
    (ain==511) ? 32'h3fb4e597 :
    (ain==512) ? 32'h3fb504f3 :
    (ain==513) ? 32'h3fb52454 :
    (ain==514) ? 32'h3fb543ba :
    (ain==515) ? 32'h3fb56326 :
    (ain==516) ? 32'h3fb58297 :
    (ain==517) ? 32'h3fb5a20e :
    (ain==518) ? 32'h3fb5c18a :
    (ain==519) ? 32'h3fb5e10c :
    (ain==520) ? 32'h3fb60093 :
    (ain==521) ? 32'h3fb62020 :
    (ain==522) ? 32'h3fb63fb2 :
    (ain==523) ? 32'h3fb65f49 :
    (ain==524) ? 32'h3fb67ee6 :
    (ain==525) ? 32'h3fb69e89 :
    (ain==526) ? 32'h3fb6be31 :
    (ain==527) ? 32'h3fb6ddde :
    (ain==528) ? 32'h3fb6fd91 :
    (ain==529) ? 32'h3fb71d4a :
    (ain==530) ? 32'h3fb73d08 :
    (ain==531) ? 32'h3fb75ccb :
    (ain==532) ? 32'h3fb77c94 :
    (ain==533) ? 32'h3fb79c63 :
    (ain==534) ? 32'h3fb7bc37 :
    (ain==535) ? 32'h3fb7dc10 :
    (ain==536) ? 32'h3fb7fbef :
    (ain==537) ? 32'h3fb81bd4 :
    (ain==538) ? 32'h3fb83bbe :
    (ain==539) ? 32'h3fb85bae :
    (ain==540) ? 32'h3fb87ba3 :
    (ain==541) ? 32'h3fb89b9d :
    (ain==542) ? 32'h3fb8bb9e :
    (ain==543) ? 32'h3fb8dba3 :
    (ain==544) ? 32'h3fb8fbaf :
    (ain==545) ? 32'h3fb91bc0 :
    (ain==546) ? 32'h3fb93bd6 :
    (ain==547) ? 32'h3fb95bf2 :
    (ain==548) ? 32'h3fb97c14 :
    (ain==549) ? 32'h3fb99c3b :
    (ain==550) ? 32'h3fb9bc68 :
    (ain==551) ? 32'h3fb9dc9a :
    (ain==552) ? 32'h3fb9fcd2 :
    (ain==553) ? 32'h3fba1d0f :
    (ain==554) ? 32'h3fba3d52 :
    (ain==555) ? 32'h3fba5d9b :
    (ain==556) ? 32'h3fba7de9 :
    (ain==557) ? 32'h3fba9e3d :
    (ain==558) ? 32'h3fbabe96 :
    (ain==559) ? 32'h3fbadef6 :
    (ain==560) ? 32'h3fbaff5a :
    (ain==561) ? 32'h3fbb1fc4 :
    (ain==562) ? 32'h3fbb4034 :
    (ain==563) ? 32'h3fbb60aa :
    (ain==564) ? 32'h3fbb8125 :
    (ain==565) ? 32'h3fbba1a6 :
    (ain==566) ? 32'h3fbbc22c :
    (ain==567) ? 32'h3fbbe2b8 :
    (ain==568) ? 32'h3fbc034a :
    (ain==569) ? 32'h3fbc23e1 :
    (ain==570) ? 32'h3fbc447e :
    (ain==571) ? 32'h3fbc6521 :
    (ain==572) ? 32'h3fbc85c9 :
    (ain==573) ? 32'h3fbca677 :
    (ain==574) ? 32'h3fbcc72b :
    (ain==575) ? 32'h3fbce7e4 :
    (ain==576) ? 32'h3fbd08a3 :
    (ain==577) ? 32'h3fbd2968 :
    (ain==578) ? 32'h3fbd4a32 :
    (ain==579) ? 32'h3fbd6b02 :
    (ain==580) ? 32'h3fbd8bd8 :
    (ain==581) ? 32'h3fbdacb3 :
    (ain==582) ? 32'h3fbdcd94 :
    (ain==583) ? 32'h3fbdee7b :
    (ain==584) ? 32'h3fbe0f68 :
    (ain==585) ? 32'h3fbe305a :
    (ain==586) ? 32'h3fbe5152 :
    (ain==587) ? 32'h3fbe724f :
    (ain==588) ? 32'h3fbe9353 :
    (ain==589) ? 32'h3fbeb45c :
    (ain==590) ? 32'h3fbed56a :
    (ain==591) ? 32'h3fbef67f :
    (ain==592) ? 32'h3fbf1799 :
    (ain==593) ? 32'h3fbf38b9 :
    (ain==594) ? 32'h3fbf59df :
    (ain==595) ? 32'h3fbf7b0a :
    (ain==596) ? 32'h3fbf9c3c :
    (ain==597) ? 32'h3fbfbd73 :
    (ain==598) ? 32'h3fbfdeaf :
    (ain==599) ? 32'h3fbffff2 :
    (ain==600) ? 32'h3fc0213a :
    (ain==601) ? 32'h3fc04288 :
    (ain==602) ? 32'h3fc063dc :
    (ain==603) ? 32'h3fc08536 :
    (ain==604) ? 32'h3fc0a695 :
    (ain==605) ? 32'h3fc0c7fa :
    (ain==606) ? 32'h3fc0e965 :
    (ain==607) ? 32'h3fc10ad6 :
    (ain==608) ? 32'h3fc12c4c :
    (ain==609) ? 32'h3fc14dc9 :
    (ain==610) ? 32'h3fc16f4b :
    (ain==611) ? 32'h3fc190d3 :
    (ain==612) ? 32'h3fc1b260 :
    (ain==613) ? 32'h3fc1d3f4 :
    (ain==614) ? 32'h3fc1f58d :
    (ain==615) ? 32'h3fc2172d :
    (ain==616) ? 32'h3fc238d2 :
    (ain==617) ? 32'h3fc25a7d :
    (ain==618) ? 32'h3fc27c2d :
    (ain==619) ? 32'h3fc29de4 :
    (ain==620) ? 32'h3fc2bfa0 :
    (ain==621) ? 32'h3fc2e162 :
    (ain==622) ? 32'h3fc3032b :
    (ain==623) ? 32'h3fc324f9 :
    (ain==624) ? 32'h3fc346cc :
    (ain==625) ? 32'h3fc368a6 :
    (ain==626) ? 32'h3fc38a86 :
    (ain==627) ? 32'h3fc3ac6b :
    (ain==628) ? 32'h3fc3ce56 :
    (ain==629) ? 32'h3fc3f047 :
    (ain==630) ? 32'h3fc4123f :
    (ain==631) ? 32'h3fc4343b :
    (ain==632) ? 32'h3fc4563e :
    (ain==633) ? 32'h3fc47847 :
    (ain==634) ? 32'h3fc49a56 :
    (ain==635) ? 32'h3fc4bc6a :
    (ain==636) ? 32'h3fc4de85 :
    (ain==637) ? 32'h3fc500a5 :
    (ain==638) ? 32'h3fc522cb :
    (ain==639) ? 32'h3fc544f7 :
    (ain==640) ? 32'h3fc5672a :
    (ain==641) ? 32'h3fc58962 :
    (ain==642) ? 32'h3fc5aba0 :
    (ain==643) ? 32'h3fc5cde3 :
    (ain==644) ? 32'h3fc5f02d :
    (ain==645) ? 32'h3fc6127d :
    (ain==646) ? 32'h3fc634d3 :
    (ain==647) ? 32'h3fc6572f :
    (ain==648) ? 32'h3fc67990 :
    (ain==649) ? 32'h3fc69bf8 :
    (ain==650) ? 32'h3fc6be65 :
    (ain==651) ? 32'h3fc6e0d9 :
    (ain==652) ? 32'h3fc70352 :
    (ain==653) ? 32'h3fc725d2 :
    (ain==654) ? 32'h3fc74857 :
    (ain==655) ? 32'h3fc76ae3 :
    (ain==656) ? 32'h3fc78d74 :
    (ain==657) ? 32'h3fc7b00c :
    (ain==658) ? 32'h3fc7d2a9 :
    (ain==659) ? 32'h3fc7f54d :
    (ain==660) ? 32'h3fc817f6 :
    (ain==661) ? 32'h3fc83aa5 :
    (ain==662) ? 32'h3fc85d5b :
    (ain==663) ? 32'h3fc88016 :
    (ain==664) ? 32'h3fc8a2d8 :
    (ain==665) ? 32'h3fc8c59f :
    (ain==666) ? 32'h3fc8e86d :
    (ain==667) ? 32'h3fc90b40 :
    (ain==668) ? 32'h3fc92e1a :
    (ain==669) ? 32'h3fc950fa :
    (ain==670) ? 32'h3fc973df :
    (ain==671) ? 32'h3fc996cb :
    (ain==672) ? 32'h3fc9b9bd :
    (ain==673) ? 32'h3fc9dcb5 :
    (ain==674) ? 32'h3fc9ffb3 :
    (ain==675) ? 32'h3fca22b7 :
    (ain==676) ? 32'h3fca45c1 :
    (ain==677) ? 32'h3fca68d1 :
    (ain==678) ? 32'h3fca8be7 :
    (ain==679) ? 32'h3fcaaf03 :
    (ain==680) ? 32'h3fcad226 :
    (ain==681) ? 32'h3fcaf54e :
    (ain==682) ? 32'h3fcb187d :
    (ain==683) ? 32'h3fcb3bb2 :
    (ain==684) ? 32'h3fcb5eec :
    (ain==685) ? 32'h3fcb822d :
    (ain==686) ? 32'h3fcba574 :
    (ain==687) ? 32'h3fcbc8c1 :
    (ain==688) ? 32'h3fcbec14 :
    (ain==689) ? 32'h3fcc0f6e :
    (ain==690) ? 32'h3fcc32cd :
    (ain==691) ? 32'h3fcc5633 :
    (ain==692) ? 32'h3fcc799f :
    (ain==693) ? 32'h3fcc9d11 :
    (ain==694) ? 32'h3fccc089 :
    (ain==695) ? 32'h3fcce407 :
    (ain==696) ? 32'h3fcd078b :
    (ain==697) ? 32'h3fcd2b16 :
    (ain==698) ? 32'h3fcd4ea6 :
    (ain==699) ? 32'h3fcd723d :
    (ain==700) ? 32'h3fcd95da :
    (ain==701) ? 32'h3fcdb97d :
    (ain==702) ? 32'h3fcddd26 :
    (ain==703) ? 32'h3fce00d6 :
    (ain==704) ? 32'h3fce248c :
    (ain==705) ? 32'h3fce4847 :
    (ain==706) ? 32'h3fce6c0a :
    (ain==707) ? 32'h3fce8fd2 :
    (ain==708) ? 32'h3fceb3a0 :
    (ain==709) ? 32'h3fced775 :
    (ain==710) ? 32'h3fcefb50 :
    (ain==711) ? 32'h3fcf1f31 :
    (ain==712) ? 32'h3fcf4318 :
    (ain==713) ? 32'h3fcf6706 :
    (ain==714) ? 32'h3fcf8afa :
    (ain==715) ? 32'h3fcfaef4 :
    (ain==716) ? 32'h3fcfd2f4 :
    (ain==717) ? 32'h3fcff6fa :
    (ain==718) ? 32'h3fd01b07 :
    (ain==719) ? 32'h3fd03f1a :
    (ain==720) ? 32'h3fd06333 :
    (ain==721) ? 32'h3fd08753 :
    (ain==722) ? 32'h3fd0ab79 :
    (ain==723) ? 32'h3fd0cfa5 :
    (ain==724) ? 32'h3fd0f3d7 :
    (ain==725) ? 32'h3fd1180f :
    (ain==726) ? 32'h3fd13c4e :
    (ain==727) ? 32'h3fd16093 :
    (ain==728) ? 32'h3fd184df :
    (ain==729) ? 32'h3fd1a931 :
    (ain==730) ? 32'h3fd1cd89 :
    (ain==731) ? 32'h3fd1f1e7 :
    (ain==732) ? 32'h3fd2164c :
    (ain==733) ? 32'h3fd23ab6 :
    (ain==734) ? 32'h3fd25f28 :
    (ain==735) ? 32'h3fd2839f :
    (ain==736) ? 32'h3fd2a81d :
    (ain==737) ? 32'h3fd2cca1 :
    (ain==738) ? 32'h3fd2f12c :
    (ain==739) ? 32'h3fd315bd :
    (ain==740) ? 32'h3fd33a54 :
    (ain==741) ? 32'h3fd35ef1 :
    (ain==742) ? 32'h3fd38395 :
    (ain==743) ? 32'h3fd3a840 :
    (ain==744) ? 32'h3fd3ccf0 :
    (ain==745) ? 32'h3fd3f1a7 :
    (ain==746) ? 32'h3fd41664 :
    (ain==747) ? 32'h3fd43b28 :
    (ain==748) ? 32'h3fd45ff2 :
    (ain==749) ? 32'h3fd484c3 :
    (ain==750) ? 32'h3fd4a999 :
    (ain==751) ? 32'h3fd4ce77 :
    (ain==752) ? 32'h3fd4f35a :
    (ain==753) ? 32'h3fd51844 :
    (ain==754) ? 32'h3fd53d35 :
    (ain==755) ? 32'h3fd5622b :
    (ain==756) ? 32'h3fd58729 :
    (ain==757) ? 32'h3fd5ac2c :
    (ain==758) ? 32'h3fd5d136 :
    (ain==759) ? 32'h3fd5f647 :
    (ain==760) ? 32'h3fd61b5d :
    (ain==761) ? 32'h3fd6407b :
    (ain==762) ? 32'h3fd6659f :
    (ain==763) ? 32'h3fd68ac9 :
    (ain==764) ? 32'h3fd6aff9 :
    (ain==765) ? 32'h3fd6d530 :
    (ain==766) ? 32'h3fd6fa6e :
    (ain==767) ? 32'h3fd71fb2 :
    (ain==768) ? 32'h3fd744fc :
    (ain==769) ? 32'h3fd76a4d :
    (ain==770) ? 32'h3fd78fa5 :
    (ain==771) ? 32'h3fd7b502 :
    (ain==772) ? 32'h3fd7da67 :
    (ain==773) ? 32'h3fd7ffd1 :
    (ain==774) ? 32'h3fd82543 :
    (ain==775) ? 32'h3fd84abb :
    (ain==776) ? 32'h3fd87039 :
    (ain==777) ? 32'h3fd895be :
    (ain==778) ? 32'h3fd8bb49 :
    (ain==779) ? 32'h3fd8e0db :
    (ain==780) ? 32'h3fd90673 :
    (ain==781) ? 32'h3fd92c12 :
    (ain==782) ? 32'h3fd951b7 :
    (ain==783) ? 32'h3fd97763 :
    (ain==784) ? 32'h3fd99d15 :
    (ain==785) ? 32'h3fd9c2ce :
    (ain==786) ? 32'h3fd9e88e :
    (ain==787) ? 32'h3fda0e54 :
    (ain==788) ? 32'h3fda3420 :
    (ain==789) ? 32'h3fda59f3 :
    (ain==790) ? 32'h3fda7fcd :
    (ain==791) ? 32'h3fdaa5ad :
    (ain==792) ? 32'h3fdacb94 :
    (ain==793) ? 32'h3fdaf181 :
    (ain==794) ? 32'h3fdb1775 :
    (ain==795) ? 32'h3fdb3d70 :
    (ain==796) ? 32'h3fdb6371 :
    (ain==797) ? 32'h3fdb8978 :
    (ain==798) ? 32'h3fdbaf87 :
    (ain==799) ? 32'h3fdbd59c :
    (ain==800) ? 32'h3fdbfbb7 :
    (ain==801) ? 32'h3fdc21d9 :
    (ain==802) ? 32'h3fdc4802 :
    (ain==803) ? 32'h3fdc6e31 :
    (ain==804) ? 32'h3fdc9467 :
    (ain==805) ? 32'h3fdcbaa4 :
    (ain==806) ? 32'h3fdce0e7 :
    (ain==807) ? 32'h3fdd0731 :
    (ain==808) ? 32'h3fdd2d81 :
    (ain==809) ? 32'h3fdd53d8 :
    (ain==810) ? 32'h3fdd7a36 :
    (ain==811) ? 32'h3fdda09a :
    (ain==812) ? 32'h3fddc705 :
    (ain==813) ? 32'h3fdded77 :
    (ain==814) ? 32'h3fde13ef :
    (ain==815) ? 32'h3fde3a6e :
    (ain==816) ? 32'h3fde60f4 :
    (ain==817) ? 32'h3fde8780 :
    (ain==818) ? 32'h3fdeae13 :
    (ain==819) ? 32'h3fded4ad :
    (ain==820) ? 32'h3fdefb4e :
    (ain==821) ? 32'h3fdf21f5 :
    (ain==822) ? 32'h3fdf48a3 :
    (ain==823) ? 32'h3fdf6f57 :
    (ain==824) ? 32'h3fdf9612 :
    (ain==825) ? 32'h3fdfbcd4 :
    (ain==826) ? 32'h3fdfe39d :
    (ain==827) ? 32'h3fe00a6c :
    (ain==828) ? 32'h3fe03143 :
    (ain==829) ? 32'h3fe0581f :
    (ain==830) ? 32'h3fe07f03 :
    (ain==831) ? 32'h3fe0a5ed :
    (ain==832) ? 32'h3fe0ccde :
    (ain==833) ? 32'h3fe0f3d6 :
    (ain==834) ? 32'h3fe11ad5 :
    (ain==835) ? 32'h3fe141da :
    (ain==836) ? 32'h3fe168e6 :
    (ain==837) ? 32'h3fe18ff9 :
    (ain==838) ? 32'h3fe1b713 :
    (ain==839) ? 32'h3fe1de33 :
    (ain==840) ? 32'h3fe2055a :
    (ain==841) ? 32'h3fe22c89 :
    (ain==842) ? 32'h3fe253bd :
    (ain==843) ? 32'h3fe27af9 :
    (ain==844) ? 32'h3fe2a23b :
    (ain==845) ? 32'h3fe2c984 :
    (ain==846) ? 32'h3fe2f0d4 :
    (ain==847) ? 32'h3fe3182b :
    (ain==848) ? 32'h3fe33f89 :
    (ain==849) ? 32'h3fe366ed :
    (ain==850) ? 32'h3fe38e59 :
    (ain==851) ? 32'h3fe3b5cb :
    (ain==852) ? 32'h3fe3dd44 :
    (ain==853) ? 32'h3fe404c4 :
    (ain==854) ? 32'h3fe42c4a :
    (ain==855) ? 32'h3fe453d8 :
    (ain==856) ? 32'h3fe47b6c :
    (ain==857) ? 32'h3fe4a307 :
    (ain==858) ? 32'h3fe4caa9 :
    (ain==859) ? 32'h3fe4f252 :
    (ain==860) ? 32'h3fe51a02 :
    (ain==861) ? 32'h3fe541b9 :
    (ain==862) ? 32'h3fe56977 :
    (ain==863) ? 32'h3fe5913b :
    (ain==864) ? 32'h3fe5b906 :
    (ain==865) ? 32'h3fe5e0d9 :
    (ain==866) ? 32'h3fe608b2 :
    (ain==867) ? 32'h3fe63092 :
    (ain==868) ? 32'h3fe65879 :
    (ain==869) ? 32'h3fe68067 :
    (ain==870) ? 32'h3fe6a85c :
    (ain==871) ? 32'h3fe6d057 :
    (ain==872) ? 32'h3fe6f85a :
    (ain==873) ? 32'h3fe72064 :
    (ain==874) ? 32'h3fe74874 :
    (ain==875) ? 32'h3fe7708c :
    (ain==876) ? 32'h3fe798aa :
    (ain==877) ? 32'h3fe7c0d0 :
    (ain==878) ? 32'h3fe7e8fc :
    (ain==879) ? 32'h3fe81130 :
    (ain==880) ? 32'h3fe8396a :
    (ain==881) ? 32'h3fe861ab :
    (ain==882) ? 32'h3fe889f3 :
    (ain==883) ? 32'h3fe8b243 :
    (ain==884) ? 32'h3fe8da99 :
    (ain==885) ? 32'h3fe902f6 :
    (ain==886) ? 32'h3fe92b5a :
    (ain==887) ? 32'h3fe953c6 :
    (ain==888) ? 32'h3fe97c38 :
    (ain==889) ? 32'h3fe9a4b1 :
    (ain==890) ? 32'h3fe9cd31 :
    (ain==891) ? 32'h3fe9f5b9 :
    (ain==892) ? 32'h3fea1e47 :
    (ain==893) ? 32'h3fea46dc :
    (ain==894) ? 32'h3fea6f79 :
    (ain==895) ? 32'h3fea981c :
    (ain==896) ? 32'h3feac0c6 :
    (ain==897) ? 32'h3feae978 :
    (ain==898) ? 32'h3feb1230 :
    (ain==899) ? 32'h3feb3af0 :
    (ain==900) ? 32'h3feb63b7 :
    (ain==901) ? 32'h3feb8c85 :
    (ain==902) ? 32'h3febb559 :
    (ain==903) ? 32'h3febde35 :
    (ain==904) ? 32'h3fec0718 :
    (ain==905) ? 32'h3fec3002 :
    (ain==906) ? 32'h3fec58f3 :
    (ain==907) ? 32'h3fec81ec :
    (ain==908) ? 32'h3fecaaeb :
    (ain==909) ? 32'h3fecd3f2 :
    (ain==910) ? 32'h3fecfcff :
    (ain==911) ? 32'h3fed2614 :
    (ain==912) ? 32'h3fed4f30 :
    (ain==913) ? 32'h3fed7853 :
    (ain==914) ? 32'h3feda17d :
    (ain==915) ? 32'h3fedcaae :
    (ain==916) ? 32'h3fedf3e6 :
    (ain==917) ? 32'h3fee1d26 :
    (ain==918) ? 32'h3fee466c :
    (ain==919) ? 32'h3fee6fba :
    (ain==920) ? 32'h3fee990f :
    (ain==921) ? 32'h3feec26b :
    (ain==922) ? 32'h3feeebcf :
    (ain==923) ? 32'h3fef1539 :
    (ain==924) ? 32'h3fef3eab :
    (ain==925) ? 32'h3fef6823 :
    (ain==926) ? 32'h3fef91a3 :
    (ain==927) ? 32'h3fefbb2b :
    (ain==928) ? 32'h3fefe4b9 :
    (ain==929) ? 32'h3ff00e4f :
    (ain==930) ? 32'h3ff037ec :
    (ain==931) ? 32'h3ff06190 :
    (ain==932) ? 32'h3ff08b3b :
    (ain==933) ? 32'h3ff0b4ed :
    (ain==934) ? 32'h3ff0dea7 :
    (ain==935) ? 32'h3ff10868 :
    (ain==936) ? 32'h3ff13230 :
    (ain==937) ? 32'h3ff15c00 :
    (ain==938) ? 32'h3ff185d6 :
    (ain==939) ? 32'h3ff1afb4 :
    (ain==940) ? 32'h3ff1d999 :
    (ain==941) ? 32'h3ff20386 :
    (ain==942) ? 32'h3ff22d79 :
    (ain==943) ? 32'h3ff25774 :
    (ain==944) ? 32'h3ff28177 :
    (ain==945) ? 32'h3ff2ab80 :
    (ain==946) ? 32'h3ff2d591 :
    (ain==947) ? 32'h3ff2ffa9 :
    (ain==948) ? 32'h3ff329c9 :
    (ain==949) ? 32'h3ff353ef :
    (ain==950) ? 32'h3ff37e1d :
    (ain==951) ? 32'h3ff3a853 :
    (ain==952) ? 32'h3ff3d28f :
    (ain==953) ? 32'h3ff3fcd3 :
    (ain==954) ? 32'h3ff4271f :
    (ain==955) ? 32'h3ff45171 :
    (ain==956) ? 32'h3ff47bcb :
    (ain==957) ? 32'h3ff4a62d :
    (ain==958) ? 32'h3ff4d095 :
    (ain==959) ? 32'h3ff4fb05 :
    (ain==960) ? 32'h3ff5257d :
    (ain==961) ? 32'h3ff54ffb :
    (ain==962) ? 32'h3ff57a81 :
    (ain==963) ? 32'h3ff5a50f :
    (ain==964) ? 32'h3ff5cfa4 :
    (ain==965) ? 32'h3ff5fa40 :
    (ain==966) ? 32'h3ff624e4 :
    (ain==967) ? 32'h3ff64f8f :
    (ain==968) ? 32'h3ff67a41 :
    (ain==969) ? 32'h3ff6a4fb :
    (ain==970) ? 32'h3ff6cfbc :
    (ain==971) ? 32'h3ff6fa85 :
    (ain==972) ? 32'h3ff72555 :
    (ain==973) ? 32'h3ff7502c :
    (ain==974) ? 32'h3ff77b0b :
    (ain==975) ? 32'h3ff7a5f1 :
    (ain==976) ? 32'h3ff7d0df :
    (ain==977) ? 32'h3ff7fbd4 :
    (ain==978) ? 32'h3ff826d1 :
    (ain==979) ? 32'h3ff851d5 :
    (ain==980) ? 32'h3ff87ce0 :
    (ain==981) ? 32'h3ff8a7f3 :
    (ain==982) ? 32'h3ff8d30e :
    (ain==983) ? 32'h3ff8fe30 :
    (ain==984) ? 32'h3ff92959 :
    (ain==985) ? 32'h3ff9548a :
    (ain==986) ? 32'h3ff97fc3 :
    (ain==987) ? 32'h3ff9ab02 :
    (ain==988) ? 32'h3ff9d64a :
    (ain==989) ? 32'h3ffa0199 :
    (ain==990) ? 32'h3ffa2cef :
    (ain==991) ? 32'h3ffa584d :
    (ain==992) ? 32'h3ffa83b2 :
    (ain==993) ? 32'h3ffaaf1f :
    (ain==994) ? 32'h3ffada94 :
    (ain==995) ? 32'h3ffb0610 :
    (ain==996) ? 32'h3ffb3193 :
    (ain==997) ? 32'h3ffb5d1e :
    (ain==998) ? 32'h3ffb88b1 :
    (ain==999) ? 32'h3ffbb44b :
    (ain==1000) ? 32'h3ffbdfed :
    (ain==1001) ? 32'h3ffc0b96 :
    (ain==1002) ? 32'h3ffc3747 :
    (ain==1003) ? 32'h3ffc6300 :
    (ain==1004) ? 32'h3ffc8ec0 :
    (ain==1005) ? 32'h3ffcba87 :
    (ain==1006) ? 32'h3ffce656 :
    (ain==1007) ? 32'h3ffd122d :
    (ain==1008) ? 32'h3ffd3e0c :
    (ain==1009) ? 32'h3ffd69f2 :
    (ain==1010) ? 32'h3ffd95df :
    (ain==1011) ? 32'h3ffdc1d4 :
    (ain==1012) ? 32'h3ffdedd1 :
    (ain==1013) ? 32'h3ffe19d6 :
    (ain==1014) ? 32'h3ffe45e2 :
    (ain==1015) ? 32'h3ffe71f5 :
    (ain==1016) ? 32'h3ffe9e11 :
    (ain==1017) ? 32'h3ffeca34 :
    (ain==1018) ? 32'h3ffef65f :
    (ain==1019) ? 32'h3fff2291 :
    (ain==1020) ? 32'h3fff4ecb :
    (ain==1021) ? 32'h3fff7b0c :
    (ain==1022) ? 32'h3fffa756 :
    (ain==1023) ? 32'h3fffd3a7 :
    0;
endmodule
