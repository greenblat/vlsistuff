
    module x16x4 #(parameter IDWID=4, parameter DWID=64, parameter EXTRAS=8, parameter WSTRB=DWID/8) ( input clk, input rst_n

    ,output [IDWID-1:0] slv0_arid
    ,output [31:0] slv0_araddr
    ,output [7:0] slv0_arlen
    ,output [2:0] slv0_arsize
    ,output [EXTRAS-1:0] slv0_arextras
    ,output [1:0] slv0_arburst
    ,output slv0_arvalid
    ,input slv0_arready
    ,input [IDWID-1:0] slv0_rid
    ,input [DWID-1:0] slv0_rdata
    ,input [1:0] slv0_rresp
    ,input slv0_rlast
    ,input slv0_rvalid
    ,output slv0_rready

    ,output [IDWID-1:0] slv0_awid
    ,output [31:0] slv0_awaddr
    ,output [7:0] slv0_awlen
    ,output [2:0] slv0_awsize
    ,output [EXTRAS-1:0] slv0_awextras
    ,output [1:0] slv0_awburst
    ,output slv0_awvalid
    ,input slv0_awready
    ,output [DWID-1:0] slv0_wdata
    ,output [WSTRB-1:0] slv0_wstrb
    ,output slv0_wlast
    ,output slv0_wvalid
    ,input slv0_wready
    ,input [IDWID-1:0] slv0_bid
    ,input [1:0] slv0_bresp
    ,input slv0_bvalid
    ,output slv0_bready

    ,output [IDWID-1:0] slv1_arid
    ,output [31:0] slv1_araddr
    ,output [7:0] slv1_arlen
    ,output [2:0] slv1_arsize
    ,output [EXTRAS-1:0] slv1_arextras
    ,output [1:0] slv1_arburst
    ,output slv1_arvalid
    ,input slv1_arready
    ,input [IDWID-1:0] slv1_rid
    ,input [DWID-1:0] slv1_rdata
    ,input [1:0] slv1_rresp
    ,input slv1_rlast
    ,input slv1_rvalid
    ,output slv1_rready

    ,output [IDWID-1:0] slv1_awid
    ,output [31:0] slv1_awaddr
    ,output [7:0] slv1_awlen
    ,output [2:0] slv1_awsize
    ,output [EXTRAS-1:0] slv1_awextras
    ,output [1:0] slv1_awburst
    ,output slv1_awvalid
    ,input slv1_awready
    ,output [DWID-1:0] slv1_wdata
    ,output [WSTRB-1:0] slv1_wstrb
    ,output slv1_wlast
    ,output slv1_wvalid
    ,input slv1_wready
    ,input [IDWID-1:0] slv1_bid
    ,input [1:0] slv1_bresp
    ,input slv1_bvalid
    ,output slv1_bready

    ,output [IDWID-1:0] slv2_arid
    ,output [31:0] slv2_araddr
    ,output [7:0] slv2_arlen
    ,output [2:0] slv2_arsize
    ,output [EXTRAS-1:0] slv2_arextras
    ,output [1:0] slv2_arburst
    ,output slv2_arvalid
    ,input slv2_arready
    ,input [IDWID-1:0] slv2_rid
    ,input [DWID-1:0] slv2_rdata
    ,input [1:0] slv2_rresp
    ,input slv2_rlast
    ,input slv2_rvalid
    ,output slv2_rready

    ,output [IDWID-1:0] slv2_awid
    ,output [31:0] slv2_awaddr
    ,output [7:0] slv2_awlen
    ,output [2:0] slv2_awsize
    ,output [EXTRAS-1:0] slv2_awextras
    ,output [1:0] slv2_awburst
    ,output slv2_awvalid
    ,input slv2_awready
    ,output [DWID-1:0] slv2_wdata
    ,output [WSTRB-1:0] slv2_wstrb
    ,output slv2_wlast
    ,output slv2_wvalid
    ,input slv2_wready
    ,input [IDWID-1:0] slv2_bid
    ,input [1:0] slv2_bresp
    ,input slv2_bvalid
    ,output slv2_bready

    ,output [IDWID-1:0] slv3_arid
    ,output [31:0] slv3_araddr
    ,output [7:0] slv3_arlen
    ,output [2:0] slv3_arsize
    ,output [EXTRAS-1:0] slv3_arextras
    ,output [1:0] slv3_arburst
    ,output slv3_arvalid
    ,input slv3_arready
    ,input [IDWID-1:0] slv3_rid
    ,input [DWID-1:0] slv3_rdata
    ,input [1:0] slv3_rresp
    ,input slv3_rlast
    ,input slv3_rvalid
    ,output slv3_rready

    ,output [IDWID-1:0] slv3_awid
    ,output [31:0] slv3_awaddr
    ,output [7:0] slv3_awlen
    ,output [2:0] slv3_awsize
    ,output [EXTRAS-1:0] slv3_awextras
    ,output [1:0] slv3_awburst
    ,output slv3_awvalid
    ,input slv3_awready
    ,output [DWID-1:0] slv3_wdata
    ,output [WSTRB-1:0] slv3_wstrb
    ,output slv3_wlast
    ,output slv3_wvalid
    ,input slv3_wready
    ,input [IDWID-1:0] slv3_bid
    ,input [1:0] slv3_bresp
    ,input slv3_bvalid
    ,output slv3_bready

    ,input [IDWID-1:0] mst0_arid
    ,input [31:0] mst0_araddr
    ,input [7:0] mst0_arlen
    ,input [2:0] mst0_arsize
    ,input [EXTRAS-1:0] mst0_arextras
    ,input [1:0] mst0_arburst
    ,input mst0_arvalid
    ,output mst0_arready
    ,output [IDWID-1:0] mst0_rid
    ,output [DWID-1:0] mst0_rdata
    ,output [1:0] mst0_rresp
    ,output mst0_rlast
    ,output mst0_rvalid
    ,input mst0_rready

    ,input [IDWID-1:0] mst0_awid
    ,input [31:0] mst0_awaddr
    ,input [7:0] mst0_awlen
    ,input [2:0] mst0_awsize
    ,input [EXTRAS-1:0] mst0_awextras
    ,input [1:0] mst0_awburst
    ,input mst0_awvalid
    ,output mst0_awready
    ,input [DWID-1:0] mst0_wdata
    ,input [WSTRB-1:0] mst0_wstrb
    ,input mst0_wlast
    ,input mst0_wvalid
    ,output mst0_wready
    ,output [IDWID-1:0] mst0_bid
    ,output [1:0] mst0_bresp
    ,output mst0_bvalid
    ,input mst0_bready

    ,input [IDWID-1:0] mst1_arid
    ,input [31:0] mst1_araddr
    ,input [7:0] mst1_arlen
    ,input [2:0] mst1_arsize
    ,input [EXTRAS-1:0] mst1_arextras
    ,input [1:0] mst1_arburst
    ,input mst1_arvalid
    ,output mst1_arready
    ,output [IDWID-1:0] mst1_rid
    ,output [DWID-1:0] mst1_rdata
    ,output [1:0] mst1_rresp
    ,output mst1_rlast
    ,output mst1_rvalid
    ,input mst1_rready

    ,input [IDWID-1:0] mst1_awid
    ,input [31:0] mst1_awaddr
    ,input [7:0] mst1_awlen
    ,input [2:0] mst1_awsize
    ,input [EXTRAS-1:0] mst1_awextras
    ,input [1:0] mst1_awburst
    ,input mst1_awvalid
    ,output mst1_awready
    ,input [DWID-1:0] mst1_wdata
    ,input [WSTRB-1:0] mst1_wstrb
    ,input mst1_wlast
    ,input mst1_wvalid
    ,output mst1_wready
    ,output [IDWID-1:0] mst1_bid
    ,output [1:0] mst1_bresp
    ,output mst1_bvalid
    ,input mst1_bready

    ,input [IDWID-1:0] mst10_arid
    ,input [31:0] mst10_araddr
    ,input [7:0] mst10_arlen
    ,input [2:0] mst10_arsize
    ,input [EXTRAS-1:0] mst10_arextras
    ,input [1:0] mst10_arburst
    ,input mst10_arvalid
    ,output mst10_arready
    ,output [IDWID-1:0] mst10_rid
    ,output [DWID-1:0] mst10_rdata
    ,output [1:0] mst10_rresp
    ,output mst10_rlast
    ,output mst10_rvalid
    ,input mst10_rready

    ,input [IDWID-1:0] mst10_awid
    ,input [31:0] mst10_awaddr
    ,input [7:0] mst10_awlen
    ,input [2:0] mst10_awsize
    ,input [EXTRAS-1:0] mst10_awextras
    ,input [1:0] mst10_awburst
    ,input mst10_awvalid
    ,output mst10_awready
    ,input [DWID-1:0] mst10_wdata
    ,input [WSTRB-1:0] mst10_wstrb
    ,input mst10_wlast
    ,input mst10_wvalid
    ,output mst10_wready
    ,output [IDWID-1:0] mst10_bid
    ,output [1:0] mst10_bresp
    ,output mst10_bvalid
    ,input mst10_bready

    ,input [IDWID-1:0] mst11_arid
    ,input [31:0] mst11_araddr
    ,input [7:0] mst11_arlen
    ,input [2:0] mst11_arsize
    ,input [EXTRAS-1:0] mst11_arextras
    ,input [1:0] mst11_arburst
    ,input mst11_arvalid
    ,output mst11_arready
    ,output [IDWID-1:0] mst11_rid
    ,output [DWID-1:0] mst11_rdata
    ,output [1:0] mst11_rresp
    ,output mst11_rlast
    ,output mst11_rvalid
    ,input mst11_rready

    ,input [IDWID-1:0] mst11_awid
    ,input [31:0] mst11_awaddr
    ,input [7:0] mst11_awlen
    ,input [2:0] mst11_awsize
    ,input [EXTRAS-1:0] mst11_awextras
    ,input [1:0] mst11_awburst
    ,input mst11_awvalid
    ,output mst11_awready
    ,input [DWID-1:0] mst11_wdata
    ,input [WSTRB-1:0] mst11_wstrb
    ,input mst11_wlast
    ,input mst11_wvalid
    ,output mst11_wready
    ,output [IDWID-1:0] mst11_bid
    ,output [1:0] mst11_bresp
    ,output mst11_bvalid
    ,input mst11_bready

    ,input [IDWID-1:0] mst12_arid
    ,input [31:0] mst12_araddr
    ,input [7:0] mst12_arlen
    ,input [2:0] mst12_arsize
    ,input [EXTRAS-1:0] mst12_arextras
    ,input [1:0] mst12_arburst
    ,input mst12_arvalid
    ,output mst12_arready
    ,output [IDWID-1:0] mst12_rid
    ,output [DWID-1:0] mst12_rdata
    ,output [1:0] mst12_rresp
    ,output mst12_rlast
    ,output mst12_rvalid
    ,input mst12_rready

    ,input [IDWID-1:0] mst12_awid
    ,input [31:0] mst12_awaddr
    ,input [7:0] mst12_awlen
    ,input [2:0] mst12_awsize
    ,input [EXTRAS-1:0] mst12_awextras
    ,input [1:0] mst12_awburst
    ,input mst12_awvalid
    ,output mst12_awready
    ,input [DWID-1:0] mst12_wdata
    ,input [WSTRB-1:0] mst12_wstrb
    ,input mst12_wlast
    ,input mst12_wvalid
    ,output mst12_wready
    ,output [IDWID-1:0] mst12_bid
    ,output [1:0] mst12_bresp
    ,output mst12_bvalid
    ,input mst12_bready

    ,input [IDWID-1:0] mst13_arid
    ,input [31:0] mst13_araddr
    ,input [7:0] mst13_arlen
    ,input [2:0] mst13_arsize
    ,input [EXTRAS-1:0] mst13_arextras
    ,input [1:0] mst13_arburst
    ,input mst13_arvalid
    ,output mst13_arready
    ,output [IDWID-1:0] mst13_rid
    ,output [DWID-1:0] mst13_rdata
    ,output [1:0] mst13_rresp
    ,output mst13_rlast
    ,output mst13_rvalid
    ,input mst13_rready

    ,input [IDWID-1:0] mst13_awid
    ,input [31:0] mst13_awaddr
    ,input [7:0] mst13_awlen
    ,input [2:0] mst13_awsize
    ,input [EXTRAS-1:0] mst13_awextras
    ,input [1:0] mst13_awburst
    ,input mst13_awvalid
    ,output mst13_awready
    ,input [DWID-1:0] mst13_wdata
    ,input [WSTRB-1:0] mst13_wstrb
    ,input mst13_wlast
    ,input mst13_wvalid
    ,output mst13_wready
    ,output [IDWID-1:0] mst13_bid
    ,output [1:0] mst13_bresp
    ,output mst13_bvalid
    ,input mst13_bready

    ,input [IDWID-1:0] mst14_arid
    ,input [31:0] mst14_araddr
    ,input [7:0] mst14_arlen
    ,input [2:0] mst14_arsize
    ,input [EXTRAS-1:0] mst14_arextras
    ,input [1:0] mst14_arburst
    ,input mst14_arvalid
    ,output mst14_arready
    ,output [IDWID-1:0] mst14_rid
    ,output [DWID-1:0] mst14_rdata
    ,output [1:0] mst14_rresp
    ,output mst14_rlast
    ,output mst14_rvalid
    ,input mst14_rready

    ,input [IDWID-1:0] mst14_awid
    ,input [31:0] mst14_awaddr
    ,input [7:0] mst14_awlen
    ,input [2:0] mst14_awsize
    ,input [EXTRAS-1:0] mst14_awextras
    ,input [1:0] mst14_awburst
    ,input mst14_awvalid
    ,output mst14_awready
    ,input [DWID-1:0] mst14_wdata
    ,input [WSTRB-1:0] mst14_wstrb
    ,input mst14_wlast
    ,input mst14_wvalid
    ,output mst14_wready
    ,output [IDWID-1:0] mst14_bid
    ,output [1:0] mst14_bresp
    ,output mst14_bvalid
    ,input mst14_bready

    ,input [IDWID-1:0] mst15_arid
    ,input [31:0] mst15_araddr
    ,input [7:0] mst15_arlen
    ,input [2:0] mst15_arsize
    ,input [EXTRAS-1:0] mst15_arextras
    ,input [1:0] mst15_arburst
    ,input mst15_arvalid
    ,output mst15_arready
    ,output [IDWID-1:0] mst15_rid
    ,output [DWID-1:0] mst15_rdata
    ,output [1:0] mst15_rresp
    ,output mst15_rlast
    ,output mst15_rvalid
    ,input mst15_rready

    ,input [IDWID-1:0] mst15_awid
    ,input [31:0] mst15_awaddr
    ,input [7:0] mst15_awlen
    ,input [2:0] mst15_awsize
    ,input [EXTRAS-1:0] mst15_awextras
    ,input [1:0] mst15_awburst
    ,input mst15_awvalid
    ,output mst15_awready
    ,input [DWID-1:0] mst15_wdata
    ,input [WSTRB-1:0] mst15_wstrb
    ,input mst15_wlast
    ,input mst15_wvalid
    ,output mst15_wready
    ,output [IDWID-1:0] mst15_bid
    ,output [1:0] mst15_bresp
    ,output mst15_bvalid
    ,input mst15_bready

    ,input [IDWID-1:0] mst2_arid
    ,input [31:0] mst2_araddr
    ,input [7:0] mst2_arlen
    ,input [2:0] mst2_arsize
    ,input [EXTRAS-1:0] mst2_arextras
    ,input [1:0] mst2_arburst
    ,input mst2_arvalid
    ,output mst2_arready
    ,output [IDWID-1:0] mst2_rid
    ,output [DWID-1:0] mst2_rdata
    ,output [1:0] mst2_rresp
    ,output mst2_rlast
    ,output mst2_rvalid
    ,input mst2_rready

    ,input [IDWID-1:0] mst2_awid
    ,input [31:0] mst2_awaddr
    ,input [7:0] mst2_awlen
    ,input [2:0] mst2_awsize
    ,input [EXTRAS-1:0] mst2_awextras
    ,input [1:0] mst2_awburst
    ,input mst2_awvalid
    ,output mst2_awready
    ,input [DWID-1:0] mst2_wdata
    ,input [WSTRB-1:0] mst2_wstrb
    ,input mst2_wlast
    ,input mst2_wvalid
    ,output mst2_wready
    ,output [IDWID-1:0] mst2_bid
    ,output [1:0] mst2_bresp
    ,output mst2_bvalid
    ,input mst2_bready

    ,input [IDWID-1:0] mst3_arid
    ,input [31:0] mst3_araddr
    ,input [7:0] mst3_arlen
    ,input [2:0] mst3_arsize
    ,input [EXTRAS-1:0] mst3_arextras
    ,input [1:0] mst3_arburst
    ,input mst3_arvalid
    ,output mst3_arready
    ,output [IDWID-1:0] mst3_rid
    ,output [DWID-1:0] mst3_rdata
    ,output [1:0] mst3_rresp
    ,output mst3_rlast
    ,output mst3_rvalid
    ,input mst3_rready

    ,input [IDWID-1:0] mst3_awid
    ,input [31:0] mst3_awaddr
    ,input [7:0] mst3_awlen
    ,input [2:0] mst3_awsize
    ,input [EXTRAS-1:0] mst3_awextras
    ,input [1:0] mst3_awburst
    ,input mst3_awvalid
    ,output mst3_awready
    ,input [DWID-1:0] mst3_wdata
    ,input [WSTRB-1:0] mst3_wstrb
    ,input mst3_wlast
    ,input mst3_wvalid
    ,output mst3_wready
    ,output [IDWID-1:0] mst3_bid
    ,output [1:0] mst3_bresp
    ,output mst3_bvalid
    ,input mst3_bready

    ,input [IDWID-1:0] mst4_arid
    ,input [31:0] mst4_araddr
    ,input [7:0] mst4_arlen
    ,input [2:0] mst4_arsize
    ,input [EXTRAS-1:0] mst4_arextras
    ,input [1:0] mst4_arburst
    ,input mst4_arvalid
    ,output mst4_arready
    ,output [IDWID-1:0] mst4_rid
    ,output [DWID-1:0] mst4_rdata
    ,output [1:0] mst4_rresp
    ,output mst4_rlast
    ,output mst4_rvalid
    ,input mst4_rready

    ,input [IDWID-1:0] mst4_awid
    ,input [31:0] mst4_awaddr
    ,input [7:0] mst4_awlen
    ,input [2:0] mst4_awsize
    ,input [EXTRAS-1:0] mst4_awextras
    ,input [1:0] mst4_awburst
    ,input mst4_awvalid
    ,output mst4_awready
    ,input [DWID-1:0] mst4_wdata
    ,input [WSTRB-1:0] mst4_wstrb
    ,input mst4_wlast
    ,input mst4_wvalid
    ,output mst4_wready
    ,output [IDWID-1:0] mst4_bid
    ,output [1:0] mst4_bresp
    ,output mst4_bvalid
    ,input mst4_bready

    ,input [IDWID-1:0] mst5_arid
    ,input [31:0] mst5_araddr
    ,input [7:0] mst5_arlen
    ,input [2:0] mst5_arsize
    ,input [EXTRAS-1:0] mst5_arextras
    ,input [1:0] mst5_arburst
    ,input mst5_arvalid
    ,output mst5_arready
    ,output [IDWID-1:0] mst5_rid
    ,output [DWID-1:0] mst5_rdata
    ,output [1:0] mst5_rresp
    ,output mst5_rlast
    ,output mst5_rvalid
    ,input mst5_rready

    ,input [IDWID-1:0] mst5_awid
    ,input [31:0] mst5_awaddr
    ,input [7:0] mst5_awlen
    ,input [2:0] mst5_awsize
    ,input [EXTRAS-1:0] mst5_awextras
    ,input [1:0] mst5_awburst
    ,input mst5_awvalid
    ,output mst5_awready
    ,input [DWID-1:0] mst5_wdata
    ,input [WSTRB-1:0] mst5_wstrb
    ,input mst5_wlast
    ,input mst5_wvalid
    ,output mst5_wready
    ,output [IDWID-1:0] mst5_bid
    ,output [1:0] mst5_bresp
    ,output mst5_bvalid
    ,input mst5_bready

    ,input [IDWID-1:0] mst6_arid
    ,input [31:0] mst6_araddr
    ,input [7:0] mst6_arlen
    ,input [2:0] mst6_arsize
    ,input [EXTRAS-1:0] mst6_arextras
    ,input [1:0] mst6_arburst
    ,input mst6_arvalid
    ,output mst6_arready
    ,output [IDWID-1:0] mst6_rid
    ,output [DWID-1:0] mst6_rdata
    ,output [1:0] mst6_rresp
    ,output mst6_rlast
    ,output mst6_rvalid
    ,input mst6_rready

    ,input [IDWID-1:0] mst6_awid
    ,input [31:0] mst6_awaddr
    ,input [7:0] mst6_awlen
    ,input [2:0] mst6_awsize
    ,input [EXTRAS-1:0] mst6_awextras
    ,input [1:0] mst6_awburst
    ,input mst6_awvalid
    ,output mst6_awready
    ,input [DWID-1:0] mst6_wdata
    ,input [WSTRB-1:0] mst6_wstrb
    ,input mst6_wlast
    ,input mst6_wvalid
    ,output mst6_wready
    ,output [IDWID-1:0] mst6_bid
    ,output [1:0] mst6_bresp
    ,output mst6_bvalid
    ,input mst6_bready

    ,input [IDWID-1:0] mst7_arid
    ,input [31:0] mst7_araddr
    ,input [7:0] mst7_arlen
    ,input [2:0] mst7_arsize
    ,input [EXTRAS-1:0] mst7_arextras
    ,input [1:0] mst7_arburst
    ,input mst7_arvalid
    ,output mst7_arready
    ,output [IDWID-1:0] mst7_rid
    ,output [DWID-1:0] mst7_rdata
    ,output [1:0] mst7_rresp
    ,output mst7_rlast
    ,output mst7_rvalid
    ,input mst7_rready

    ,input [IDWID-1:0] mst7_awid
    ,input [31:0] mst7_awaddr
    ,input [7:0] mst7_awlen
    ,input [2:0] mst7_awsize
    ,input [EXTRAS-1:0] mst7_awextras
    ,input [1:0] mst7_awburst
    ,input mst7_awvalid
    ,output mst7_awready
    ,input [DWID-1:0] mst7_wdata
    ,input [WSTRB-1:0] mst7_wstrb
    ,input mst7_wlast
    ,input mst7_wvalid
    ,output mst7_wready
    ,output [IDWID-1:0] mst7_bid
    ,output [1:0] mst7_bresp
    ,output mst7_bvalid
    ,input mst7_bready

    ,input [IDWID-1:0] mst8_arid
    ,input [31:0] mst8_araddr
    ,input [7:0] mst8_arlen
    ,input [2:0] mst8_arsize
    ,input [EXTRAS-1:0] mst8_arextras
    ,input [1:0] mst8_arburst
    ,input mst8_arvalid
    ,output mst8_arready
    ,output [IDWID-1:0] mst8_rid
    ,output [DWID-1:0] mst8_rdata
    ,output [1:0] mst8_rresp
    ,output mst8_rlast
    ,output mst8_rvalid
    ,input mst8_rready

    ,input [IDWID-1:0] mst8_awid
    ,input [31:0] mst8_awaddr
    ,input [7:0] mst8_awlen
    ,input [2:0] mst8_awsize
    ,input [EXTRAS-1:0] mst8_awextras
    ,input [1:0] mst8_awburst
    ,input mst8_awvalid
    ,output mst8_awready
    ,input [DWID-1:0] mst8_wdata
    ,input [WSTRB-1:0] mst8_wstrb
    ,input mst8_wlast
    ,input mst8_wvalid
    ,output mst8_wready
    ,output [IDWID-1:0] mst8_bid
    ,output [1:0] mst8_bresp
    ,output mst8_bvalid
    ,input mst8_bready

    ,input [IDWID-1:0] mst9_arid
    ,input [31:0] mst9_araddr
    ,input [7:0] mst9_arlen
    ,input [2:0] mst9_arsize
    ,input [EXTRAS-1:0] mst9_arextras
    ,input [1:0] mst9_arburst
    ,input mst9_arvalid
    ,output mst9_arready
    ,output [IDWID-1:0] mst9_rid
    ,output [DWID-1:0] mst9_rdata
    ,output [1:0] mst9_rresp
    ,output mst9_rlast
    ,output mst9_rvalid
    ,input mst9_rready

    ,input [IDWID-1:0] mst9_awid
    ,input [31:0] mst9_awaddr
    ,input [7:0] mst9_awlen
    ,input [2:0] mst9_awsize
    ,input [EXTRAS-1:0] mst9_awextras
    ,input [1:0] mst9_awburst
    ,input mst9_awvalid
    ,output mst9_awready
    ,input [DWID-1:0] mst9_wdata
    ,input [WSTRB-1:0] mst9_wstrb
    ,input mst9_wlast
    ,input mst9_wvalid
    ,output mst9_wready
    ,output [IDWID-1:0] mst9_bid
    ,output [1:0] mst9_bresp
    ,output mst9_bvalid
    ,input mst9_bready
);

wire [IDWID-1:0] merger0_merger4_arid ;
wire [31:0] merger0_merger4_araddr ;
wire [7:0] merger0_merger4_arlen ;
wire [2:0] merger0_merger4_arsize ;
wire [EXTRAS-1:0] merger0_merger4_arextras ;
wire [1:0] merger0_merger4_arburst ;
wire merger0_merger4_arvalid ;
wire merger0_merger4_arready ;
wire [IDWID-1:0] merger0_merger4_rid ;
wire [DWID-1:0] merger0_merger4_rdata ;
wire [1:0] merger0_merger4_rresp ;
wire merger0_merger4_rlast ;
wire merger0_merger4_rvalid ;
wire merger0_merger4_rready ;

wire [IDWID-1:0] merger0_merger4_awid ;
wire [31:0] merger0_merger4_awaddr ;
wire [7:0] merger0_merger4_awlen ;
wire [2:0] merger0_merger4_awsize ;
wire [EXTRAS-1:0] merger0_merger4_awextras ;
wire [1:0] merger0_merger4_awburst ;
wire merger0_merger4_awvalid ;
wire merger0_merger4_awready ;
wire [DWID-1:0] merger0_merger4_wdata ;
wire [WSTRB-1:0] merger0_merger4_wstrb ;
wire merger0_merger4_wlast ;
wire merger0_merger4_wvalid ;
wire merger0_merger4_wready ;
wire [IDWID-1:0] merger0_merger4_bid ;
wire [1:0] merger0_merger4_bresp ;
wire merger0_merger4_bvalid ;
wire merger0_merger4_bready ;


axi_4_merger merger0 (
     .clk(clk),.rst_n(rst_n)
    ,.araddr(merger0_merger4_araddr[31:0])
    ,.arburst(merger0_merger4_arburst[1:0])
    ,.arextras(merger0_merger4_arextras[(EXTRAS - 1):0])
    ,.arid(merger0_merger4_arid)
    ,.arlen(merger0_merger4_arlen)
    ,.arsize(merger0_merger4_arsize)
    ,.arready(merger0_merger4_arready)
    ,.arvalid(merger0_merger4_arvalid)
    ,.awaddr(merger0_merger4_awaddr[31:0])
    ,.awburst(merger0_merger4_awburst[1:0])
    ,.awextras(merger0_merger4_awextras[(EXTRAS - 1):0])
    ,.awid(merger0_merger4_awid)
    ,.awlen(merger0_merger4_awlen)
    ,.awsize(merger0_merger4_awsize)
    ,.awready(merger0_merger4_awready)
    ,.awvalid(merger0_merger4_awvalid)
    ,.bid(merger0_merger4_bid[(IDWID - 1):0])
    ,.bready(merger0_merger4_bready)
    ,.bresp(merger0_merger4_bresp[1:0])
    ,.bvalid(merger0_merger4_bvalid)
    ,.rid(merger0_merger4_rid[(IDWID - 1):0])
    ,.rlast(merger0_merger4_rlast)
    ,.rready(merger0_merger4_rready)
    ,.rresp(merger0_merger4_rresp[1:0])
    ,.rvalid(merger0_merger4_rvalid)
    ,.rdata(merger0_merger4_rdata[(DWID - 1):0])
    ,.wdata(merger0_merger4_wdata[(DWID - 1):0])
    ,.wlast(merger0_merger4_wlast)
    ,.wready(merger0_merger4_wready)
    ,.wstrb(merger0_merger4_wstrb[(WSTRB - 1):0])
    ,.wvalid(merger0_merger4_wvalid)


    ,.a_araddr(mst0_araddr[31:0])
    ,.a_arburst(mst0_arburst[1:0])
    ,.a_arextras(mst0_arextras[(EXTRAS - 1):0])
    ,.a_arid(mst0_arid)
    ,.a_arlen(mst0_arlen)
    ,.a_arsize(mst0_arsize)
    ,.a_arready(mst0_arready)
    ,.a_arvalid(mst0_arvalid)
    ,.a_awaddr(mst0_awaddr[31:0])
    ,.a_awburst(mst0_awburst[1:0])
    ,.a_awextras(mst0_awextras[(EXTRAS - 1):0])
    ,.a_awid(mst0_awid)
    ,.a_awlen(mst0_awlen)
    ,.a_awsize(mst0_awsize)
    ,.a_awready(mst0_awready)
    ,.a_awvalid(mst0_awvalid)
    ,.a_bid(mst0_bid[(IDWID - 1):0])
    ,.a_bready(mst0_bready)
    ,.a_bresp(mst0_bresp[1:0])
    ,.a_bvalid(mst0_bvalid)
    ,.a_rdata(mst0_rdata[(DWID - 1):0])
    ,.a_rid(mst0_rid[(IDWID - 1):0])
    ,.a_rlast(mst0_rlast)
    ,.a_rready(mst0_rready)
    ,.a_rresp(mst0_rresp[1:0])
    ,.a_rvalid(mst0_rvalid)
    ,.a_wdata(mst0_wdata[(DWID - 1):0])
    ,.a_wlast(mst0_wlast)
    ,.a_wready(mst0_wready)
    ,.a_wstrb(mst0_wstrb[(WSTRB - 1):0])
    ,.a_wvalid(mst0_wvalid)

    ,.b_araddr(mst1_araddr[31:0])
    ,.b_arburst(mst1_arburst[1:0])
    ,.b_arextras(mst1_arextras[(EXTRAS - 1):0])
    ,.b_arid(mst1_arid)
    ,.b_arlen(mst1_arlen)
    ,.b_arsize(mst1_arsize)
    ,.b_arready(mst1_arready)
    ,.b_arvalid(mst1_arvalid)
    ,.b_awaddr(mst1_awaddr[31:0])
    ,.b_awburst(mst1_awburst[1:0])
    ,.b_awextras(mst1_awextras[(EXTRAS - 1):0])
    ,.b_awid(mst1_awid)
    ,.b_awlen(mst1_awlen)
    ,.b_awsize(mst1_awsize)
    ,.b_awready(mst1_awready)
    ,.b_awvalid(mst1_awvalid)
    ,.b_bid(mst1_bid[(IDWID - 1):0])
    ,.b_bready(mst1_bready)
    ,.b_bresp(mst1_bresp[1:0])
    ,.b_bvalid(mst1_bvalid)
    ,.b_rdata(mst1_rdata[(DWID - 1):0])
    ,.b_rid(mst1_rid[(IDWID - 1):0])
    ,.b_rlast(mst1_rlast)
    ,.b_rready(mst1_rready)
    ,.b_rresp(mst1_rresp[1:0])
    ,.b_rvalid(mst1_rvalid)
    ,.b_wdata(mst1_wdata[(DWID - 1):0])
    ,.b_wlast(mst1_wlast)
    ,.b_wready(mst1_wready)
    ,.b_wstrb(mst1_wstrb[(WSTRB - 1):0])
    ,.b_wvalid(mst1_wvalid)

    ,.c_araddr(mst2_araddr[31:0])
    ,.c_arburst(mst2_arburst[1:0])
    ,.c_arextras(mst2_arextras[(EXTRAS - 1):0])
    ,.c_arid(mst2_arid)
    ,.c_arlen(mst2_arlen)
    ,.c_arsize(mst2_arsize)
    ,.c_arready(mst2_arready)
    ,.c_arvalid(mst2_arvalid)
    ,.c_awaddr(mst2_awaddr[31:0])
    ,.c_awburst(mst2_awburst[1:0])
    ,.c_awextras(mst2_awextras[(EXTRAS - 1):0])
    ,.c_awid(mst2_awid)
    ,.c_awlen(mst2_awlen)
    ,.c_awsize(mst2_awsize)
    ,.c_awready(mst2_awready)
    ,.c_awvalid(mst2_awvalid)
    ,.c_bid(mst2_bid[(IDWID - 1):0])
    ,.c_bready(mst2_bready)
    ,.c_bresp(mst2_bresp[1:0])
    ,.c_bvalid(mst2_bvalid)
    ,.c_rdata(mst2_rdata[(DWID - 1):0])
    ,.c_rid(mst2_rid[(IDWID - 1):0])
    ,.c_rlast(mst2_rlast)
    ,.c_rready(mst2_rready)
    ,.c_rresp(mst2_rresp[1:0])
    ,.c_rvalid(mst2_rvalid)
    ,.c_wdata(mst2_wdata[(DWID - 1):0])
    ,.c_wlast(mst2_wlast)
    ,.c_wready(mst2_wready)
    ,.c_wstrb(mst2_wstrb[(WSTRB - 1):0])
    ,.c_wvalid(mst2_wvalid)

    ,.d_araddr(mst3_araddr[31:0])
    ,.d_arburst(mst3_arburst[1:0])
    ,.d_arextras(mst3_arextras[(EXTRAS - 1):0])
    ,.d_arid(mst3_arid)
    ,.d_arlen(mst3_arlen)
    ,.d_arsize(mst3_arsize)
    ,.d_arready(mst3_arready)
    ,.d_arvalid(mst3_arvalid)
    ,.d_awaddr(mst3_awaddr[31:0])
    ,.d_awburst(mst3_awburst[1:0])
    ,.d_awextras(mst3_awextras[(EXTRAS - 1):0])
    ,.d_awid(mst3_awid)
    ,.d_awlen(mst3_awlen)
    ,.d_awsize(mst3_awsize)
    ,.d_awready(mst3_awready)
    ,.d_awvalid(mst3_awvalid)
    ,.d_bid(mst3_bid[(IDWID - 1):0])
    ,.d_bready(mst3_bready)
    ,.d_bresp(mst3_bresp[1:0])
    ,.d_bvalid(mst3_bvalid)
    ,.d_rdata(mst3_rdata[(DWID - 1):0])
    ,.d_rid(mst3_rid[(IDWID - 1):0])
    ,.d_rlast(mst3_rlast)
    ,.d_rready(mst3_rready)
    ,.d_rresp(mst3_rresp[1:0])
    ,.d_rvalid(mst3_rvalid)
    ,.d_wdata(mst3_wdata[(DWID - 1):0])
    ,.d_wlast(mst3_wlast)
    ,.d_wready(mst3_wready)
    ,.d_wstrb(mst3_wstrb[(WSTRB - 1):0])
    ,.d_wvalid(mst3_wvalid)
);


wire [IDWID-1:0] merger1_merger4_arid ;
wire [31:0] merger1_merger4_araddr ;
wire [7:0] merger1_merger4_arlen ;
wire [2:0] merger1_merger4_arsize ;
wire [EXTRAS-1:0] merger1_merger4_arextras ;
wire [1:0] merger1_merger4_arburst ;
wire merger1_merger4_arvalid ;
wire merger1_merger4_arready ;
wire [IDWID-1:0] merger1_merger4_rid ;
wire [DWID-1:0] merger1_merger4_rdata ;
wire [1:0] merger1_merger4_rresp ;
wire merger1_merger4_rlast ;
wire merger1_merger4_rvalid ;
wire merger1_merger4_rready ;

wire [IDWID-1:0] merger1_merger4_awid ;
wire [31:0] merger1_merger4_awaddr ;
wire [7:0] merger1_merger4_awlen ;
wire [2:0] merger1_merger4_awsize ;
wire [EXTRAS-1:0] merger1_merger4_awextras ;
wire [1:0] merger1_merger4_awburst ;
wire merger1_merger4_awvalid ;
wire merger1_merger4_awready ;
wire [DWID-1:0] merger1_merger4_wdata ;
wire [WSTRB-1:0] merger1_merger4_wstrb ;
wire merger1_merger4_wlast ;
wire merger1_merger4_wvalid ;
wire merger1_merger4_wready ;
wire [IDWID-1:0] merger1_merger4_bid ;
wire [1:0] merger1_merger4_bresp ;
wire merger1_merger4_bvalid ;
wire merger1_merger4_bready ;


axi_4_merger merger1 (
     .clk(clk),.rst_n(rst_n)
    ,.araddr(merger1_merger4_araddr[31:0])
    ,.arburst(merger1_merger4_arburst[1:0])
    ,.arextras(merger1_merger4_arextras[(EXTRAS - 1):0])
    ,.arid(merger1_merger4_arid)
    ,.arlen(merger1_merger4_arlen)
    ,.arsize(merger1_merger4_arsize)
    ,.arready(merger1_merger4_arready)
    ,.arvalid(merger1_merger4_arvalid)
    ,.awaddr(merger1_merger4_awaddr[31:0])
    ,.awburst(merger1_merger4_awburst[1:0])
    ,.awextras(merger1_merger4_awextras[(EXTRAS - 1):0])
    ,.awid(merger1_merger4_awid)
    ,.awlen(merger1_merger4_awlen)
    ,.awsize(merger1_merger4_awsize)
    ,.awready(merger1_merger4_awready)
    ,.awvalid(merger1_merger4_awvalid)
    ,.bid(merger1_merger4_bid[(IDWID - 1):0])
    ,.bready(merger1_merger4_bready)
    ,.bresp(merger1_merger4_bresp[1:0])
    ,.bvalid(merger1_merger4_bvalid)
    ,.rid(merger1_merger4_rid[(IDWID - 1):0])
    ,.rlast(merger1_merger4_rlast)
    ,.rready(merger1_merger4_rready)
    ,.rresp(merger1_merger4_rresp[1:0])
    ,.rvalid(merger1_merger4_rvalid)
    ,.rdata(merger1_merger4_rdata[(DWID - 1):0])
    ,.wdata(merger1_merger4_wdata[(DWID - 1):0])
    ,.wlast(merger1_merger4_wlast)
    ,.wready(merger1_merger4_wready)
    ,.wstrb(merger1_merger4_wstrb[(WSTRB - 1):0])
    ,.wvalid(merger1_merger4_wvalid)


    ,.a_araddr(mst4_araddr[31:0])
    ,.a_arburst(mst4_arburst[1:0])
    ,.a_arextras(mst4_arextras[(EXTRAS - 1):0])
    ,.a_arid(mst4_arid)
    ,.a_arlen(mst4_arlen)
    ,.a_arsize(mst4_arsize)
    ,.a_arready(mst4_arready)
    ,.a_arvalid(mst4_arvalid)
    ,.a_awaddr(mst4_awaddr[31:0])
    ,.a_awburst(mst4_awburst[1:0])
    ,.a_awextras(mst4_awextras[(EXTRAS - 1):0])
    ,.a_awid(mst4_awid)
    ,.a_awlen(mst4_awlen)
    ,.a_awsize(mst4_awsize)
    ,.a_awready(mst4_awready)
    ,.a_awvalid(mst4_awvalid)
    ,.a_bid(mst4_bid[(IDWID - 1):0])
    ,.a_bready(mst4_bready)
    ,.a_bresp(mst4_bresp[1:0])
    ,.a_bvalid(mst4_bvalid)
    ,.a_rdata(mst4_rdata[(DWID - 1):0])
    ,.a_rid(mst4_rid[(IDWID - 1):0])
    ,.a_rlast(mst4_rlast)
    ,.a_rready(mst4_rready)
    ,.a_rresp(mst4_rresp[1:0])
    ,.a_rvalid(mst4_rvalid)
    ,.a_wdata(mst4_wdata[(DWID - 1):0])
    ,.a_wlast(mst4_wlast)
    ,.a_wready(mst4_wready)
    ,.a_wstrb(mst4_wstrb[(WSTRB - 1):0])
    ,.a_wvalid(mst4_wvalid)

    ,.b_araddr(mst5_araddr[31:0])
    ,.b_arburst(mst5_arburst[1:0])
    ,.b_arextras(mst5_arextras[(EXTRAS - 1):0])
    ,.b_arid(mst5_arid)
    ,.b_arlen(mst5_arlen)
    ,.b_arsize(mst5_arsize)
    ,.b_arready(mst5_arready)
    ,.b_arvalid(mst5_arvalid)
    ,.b_awaddr(mst5_awaddr[31:0])
    ,.b_awburst(mst5_awburst[1:0])
    ,.b_awextras(mst5_awextras[(EXTRAS - 1):0])
    ,.b_awid(mst5_awid)
    ,.b_awlen(mst5_awlen)
    ,.b_awsize(mst5_awsize)
    ,.b_awready(mst5_awready)
    ,.b_awvalid(mst5_awvalid)
    ,.b_bid(mst5_bid[(IDWID - 1):0])
    ,.b_bready(mst5_bready)
    ,.b_bresp(mst5_bresp[1:0])
    ,.b_bvalid(mst5_bvalid)
    ,.b_rdata(mst5_rdata[(DWID - 1):0])
    ,.b_rid(mst5_rid[(IDWID - 1):0])
    ,.b_rlast(mst5_rlast)
    ,.b_rready(mst5_rready)
    ,.b_rresp(mst5_rresp[1:0])
    ,.b_rvalid(mst5_rvalid)
    ,.b_wdata(mst5_wdata[(DWID - 1):0])
    ,.b_wlast(mst5_wlast)
    ,.b_wready(mst5_wready)
    ,.b_wstrb(mst5_wstrb[(WSTRB - 1):0])
    ,.b_wvalid(mst5_wvalid)

    ,.c_araddr(mst6_araddr[31:0])
    ,.c_arburst(mst6_arburst[1:0])
    ,.c_arextras(mst6_arextras[(EXTRAS - 1):0])
    ,.c_arid(mst6_arid)
    ,.c_arlen(mst6_arlen)
    ,.c_arsize(mst6_arsize)
    ,.c_arready(mst6_arready)
    ,.c_arvalid(mst6_arvalid)
    ,.c_awaddr(mst6_awaddr[31:0])
    ,.c_awburst(mst6_awburst[1:0])
    ,.c_awextras(mst6_awextras[(EXTRAS - 1):0])
    ,.c_awid(mst6_awid)
    ,.c_awlen(mst6_awlen)
    ,.c_awsize(mst6_awsize)
    ,.c_awready(mst6_awready)
    ,.c_awvalid(mst6_awvalid)
    ,.c_bid(mst6_bid[(IDWID - 1):0])
    ,.c_bready(mst6_bready)
    ,.c_bresp(mst6_bresp[1:0])
    ,.c_bvalid(mst6_bvalid)
    ,.c_rdata(mst6_rdata[(DWID - 1):0])
    ,.c_rid(mst6_rid[(IDWID - 1):0])
    ,.c_rlast(mst6_rlast)
    ,.c_rready(mst6_rready)
    ,.c_rresp(mst6_rresp[1:0])
    ,.c_rvalid(mst6_rvalid)
    ,.c_wdata(mst6_wdata[(DWID - 1):0])
    ,.c_wlast(mst6_wlast)
    ,.c_wready(mst6_wready)
    ,.c_wstrb(mst6_wstrb[(WSTRB - 1):0])
    ,.c_wvalid(mst6_wvalid)

    ,.d_araddr(mst7_araddr[31:0])
    ,.d_arburst(mst7_arburst[1:0])
    ,.d_arextras(mst7_arextras[(EXTRAS - 1):0])
    ,.d_arid(mst7_arid)
    ,.d_arlen(mst7_arlen)
    ,.d_arsize(mst7_arsize)
    ,.d_arready(mst7_arready)
    ,.d_arvalid(mst7_arvalid)
    ,.d_awaddr(mst7_awaddr[31:0])
    ,.d_awburst(mst7_awburst[1:0])
    ,.d_awextras(mst7_awextras[(EXTRAS - 1):0])
    ,.d_awid(mst7_awid)
    ,.d_awlen(mst7_awlen)
    ,.d_awsize(mst7_awsize)
    ,.d_awready(mst7_awready)
    ,.d_awvalid(mst7_awvalid)
    ,.d_bid(mst7_bid[(IDWID - 1):0])
    ,.d_bready(mst7_bready)
    ,.d_bresp(mst7_bresp[1:0])
    ,.d_bvalid(mst7_bvalid)
    ,.d_rdata(mst7_rdata[(DWID - 1):0])
    ,.d_rid(mst7_rid[(IDWID - 1):0])
    ,.d_rlast(mst7_rlast)
    ,.d_rready(mst7_rready)
    ,.d_rresp(mst7_rresp[1:0])
    ,.d_rvalid(mst7_rvalid)
    ,.d_wdata(mst7_wdata[(DWID - 1):0])
    ,.d_wlast(mst7_wlast)
    ,.d_wready(mst7_wready)
    ,.d_wstrb(mst7_wstrb[(WSTRB - 1):0])
    ,.d_wvalid(mst7_wvalid)
);


wire [IDWID-1:0] merger2_merger4_arid ;
wire [31:0] merger2_merger4_araddr ;
wire [7:0] merger2_merger4_arlen ;
wire [2:0] merger2_merger4_arsize ;
wire [EXTRAS-1:0] merger2_merger4_arextras ;
wire [1:0] merger2_merger4_arburst ;
wire merger2_merger4_arvalid ;
wire merger2_merger4_arready ;
wire [IDWID-1:0] merger2_merger4_rid ;
wire [DWID-1:0] merger2_merger4_rdata ;
wire [1:0] merger2_merger4_rresp ;
wire merger2_merger4_rlast ;
wire merger2_merger4_rvalid ;
wire merger2_merger4_rready ;

wire [IDWID-1:0] merger2_merger4_awid ;
wire [31:0] merger2_merger4_awaddr ;
wire [7:0] merger2_merger4_awlen ;
wire [2:0] merger2_merger4_awsize ;
wire [EXTRAS-1:0] merger2_merger4_awextras ;
wire [1:0] merger2_merger4_awburst ;
wire merger2_merger4_awvalid ;
wire merger2_merger4_awready ;
wire [DWID-1:0] merger2_merger4_wdata ;
wire [WSTRB-1:0] merger2_merger4_wstrb ;
wire merger2_merger4_wlast ;
wire merger2_merger4_wvalid ;
wire merger2_merger4_wready ;
wire [IDWID-1:0] merger2_merger4_bid ;
wire [1:0] merger2_merger4_bresp ;
wire merger2_merger4_bvalid ;
wire merger2_merger4_bready ;


axi_4_merger merger2 (
     .clk(clk),.rst_n(rst_n)
    ,.araddr(merger2_merger4_araddr[31:0])
    ,.arburst(merger2_merger4_arburst[1:0])
    ,.arextras(merger2_merger4_arextras[(EXTRAS - 1):0])
    ,.arid(merger2_merger4_arid)
    ,.arlen(merger2_merger4_arlen)
    ,.arsize(merger2_merger4_arsize)
    ,.arready(merger2_merger4_arready)
    ,.arvalid(merger2_merger4_arvalid)
    ,.awaddr(merger2_merger4_awaddr[31:0])
    ,.awburst(merger2_merger4_awburst[1:0])
    ,.awextras(merger2_merger4_awextras[(EXTRAS - 1):0])
    ,.awid(merger2_merger4_awid)
    ,.awlen(merger2_merger4_awlen)
    ,.awsize(merger2_merger4_awsize)
    ,.awready(merger2_merger4_awready)
    ,.awvalid(merger2_merger4_awvalid)
    ,.bid(merger2_merger4_bid[(IDWID - 1):0])
    ,.bready(merger2_merger4_bready)
    ,.bresp(merger2_merger4_bresp[1:0])
    ,.bvalid(merger2_merger4_bvalid)
    ,.rid(merger2_merger4_rid[(IDWID - 1):0])
    ,.rlast(merger2_merger4_rlast)
    ,.rready(merger2_merger4_rready)
    ,.rresp(merger2_merger4_rresp[1:0])
    ,.rvalid(merger2_merger4_rvalid)
    ,.rdata(merger2_merger4_rdata[(DWID - 1):0])
    ,.wdata(merger2_merger4_wdata[(DWID - 1):0])
    ,.wlast(merger2_merger4_wlast)
    ,.wready(merger2_merger4_wready)
    ,.wstrb(merger2_merger4_wstrb[(WSTRB - 1):0])
    ,.wvalid(merger2_merger4_wvalid)


    ,.a_araddr(mst8_araddr[31:0])
    ,.a_arburst(mst8_arburst[1:0])
    ,.a_arextras(mst8_arextras[(EXTRAS - 1):0])
    ,.a_arid(mst8_arid)
    ,.a_arlen(mst8_arlen)
    ,.a_arsize(mst8_arsize)
    ,.a_arready(mst8_arready)
    ,.a_arvalid(mst8_arvalid)
    ,.a_awaddr(mst8_awaddr[31:0])
    ,.a_awburst(mst8_awburst[1:0])
    ,.a_awextras(mst8_awextras[(EXTRAS - 1):0])
    ,.a_awid(mst8_awid)
    ,.a_awlen(mst8_awlen)
    ,.a_awsize(mst8_awsize)
    ,.a_awready(mst8_awready)
    ,.a_awvalid(mst8_awvalid)
    ,.a_bid(mst8_bid[(IDWID - 1):0])
    ,.a_bready(mst8_bready)
    ,.a_bresp(mst8_bresp[1:0])
    ,.a_bvalid(mst8_bvalid)
    ,.a_rdata(mst8_rdata[(DWID - 1):0])
    ,.a_rid(mst8_rid[(IDWID - 1):0])
    ,.a_rlast(mst8_rlast)
    ,.a_rready(mst8_rready)
    ,.a_rresp(mst8_rresp[1:0])
    ,.a_rvalid(mst8_rvalid)
    ,.a_wdata(mst8_wdata[(DWID - 1):0])
    ,.a_wlast(mst8_wlast)
    ,.a_wready(mst8_wready)
    ,.a_wstrb(mst8_wstrb[(WSTRB - 1):0])
    ,.a_wvalid(mst8_wvalid)

    ,.b_araddr(mst9_araddr[31:0])
    ,.b_arburst(mst9_arburst[1:0])
    ,.b_arextras(mst9_arextras[(EXTRAS - 1):0])
    ,.b_arid(mst9_arid)
    ,.b_arlen(mst9_arlen)
    ,.b_arsize(mst9_arsize)
    ,.b_arready(mst9_arready)
    ,.b_arvalid(mst9_arvalid)
    ,.b_awaddr(mst9_awaddr[31:0])
    ,.b_awburst(mst9_awburst[1:0])
    ,.b_awextras(mst9_awextras[(EXTRAS - 1):0])
    ,.b_awid(mst9_awid)
    ,.b_awlen(mst9_awlen)
    ,.b_awsize(mst9_awsize)
    ,.b_awready(mst9_awready)
    ,.b_awvalid(mst9_awvalid)
    ,.b_bid(mst9_bid[(IDWID - 1):0])
    ,.b_bready(mst9_bready)
    ,.b_bresp(mst9_bresp[1:0])
    ,.b_bvalid(mst9_bvalid)
    ,.b_rdata(mst9_rdata[(DWID - 1):0])
    ,.b_rid(mst9_rid[(IDWID - 1):0])
    ,.b_rlast(mst9_rlast)
    ,.b_rready(mst9_rready)
    ,.b_rresp(mst9_rresp[1:0])
    ,.b_rvalid(mst9_rvalid)
    ,.b_wdata(mst9_wdata[(DWID - 1):0])
    ,.b_wlast(mst9_wlast)
    ,.b_wready(mst9_wready)
    ,.b_wstrb(mst9_wstrb[(WSTRB - 1):0])
    ,.b_wvalid(mst9_wvalid)

    ,.c_araddr(mst10_araddr[31:0])
    ,.c_arburst(mst10_arburst[1:0])
    ,.c_arextras(mst10_arextras[(EXTRAS - 1):0])
    ,.c_arid(mst10_arid)
    ,.c_arlen(mst10_arlen)
    ,.c_arsize(mst10_arsize)
    ,.c_arready(mst10_arready)
    ,.c_arvalid(mst10_arvalid)
    ,.c_awaddr(mst10_awaddr[31:0])
    ,.c_awburst(mst10_awburst[1:0])
    ,.c_awextras(mst10_awextras[(EXTRAS - 1):0])
    ,.c_awid(mst10_awid)
    ,.c_awlen(mst10_awlen)
    ,.c_awsize(mst10_awsize)
    ,.c_awready(mst10_awready)
    ,.c_awvalid(mst10_awvalid)
    ,.c_bid(mst10_bid[(IDWID - 1):0])
    ,.c_bready(mst10_bready)
    ,.c_bresp(mst10_bresp[1:0])
    ,.c_bvalid(mst10_bvalid)
    ,.c_rdata(mst10_rdata[(DWID - 1):0])
    ,.c_rid(mst10_rid[(IDWID - 1):0])
    ,.c_rlast(mst10_rlast)
    ,.c_rready(mst10_rready)
    ,.c_rresp(mst10_rresp[1:0])
    ,.c_rvalid(mst10_rvalid)
    ,.c_wdata(mst10_wdata[(DWID - 1):0])
    ,.c_wlast(mst10_wlast)
    ,.c_wready(mst10_wready)
    ,.c_wstrb(mst10_wstrb[(WSTRB - 1):0])
    ,.c_wvalid(mst10_wvalid)

    ,.d_araddr(mst11_araddr[31:0])
    ,.d_arburst(mst11_arburst[1:0])
    ,.d_arextras(mst11_arextras[(EXTRAS - 1):0])
    ,.d_arid(mst11_arid)
    ,.d_arlen(mst11_arlen)
    ,.d_arsize(mst11_arsize)
    ,.d_arready(mst11_arready)
    ,.d_arvalid(mst11_arvalid)
    ,.d_awaddr(mst11_awaddr[31:0])
    ,.d_awburst(mst11_awburst[1:0])
    ,.d_awextras(mst11_awextras[(EXTRAS - 1):0])
    ,.d_awid(mst11_awid)
    ,.d_awlen(mst11_awlen)
    ,.d_awsize(mst11_awsize)
    ,.d_awready(mst11_awready)
    ,.d_awvalid(mst11_awvalid)
    ,.d_bid(mst11_bid[(IDWID - 1):0])
    ,.d_bready(mst11_bready)
    ,.d_bresp(mst11_bresp[1:0])
    ,.d_bvalid(mst11_bvalid)
    ,.d_rdata(mst11_rdata[(DWID - 1):0])
    ,.d_rid(mst11_rid[(IDWID - 1):0])
    ,.d_rlast(mst11_rlast)
    ,.d_rready(mst11_rready)
    ,.d_rresp(mst11_rresp[1:0])
    ,.d_rvalid(mst11_rvalid)
    ,.d_wdata(mst11_wdata[(DWID - 1):0])
    ,.d_wlast(mst11_wlast)
    ,.d_wready(mst11_wready)
    ,.d_wstrb(mst11_wstrb[(WSTRB - 1):0])
    ,.d_wvalid(mst11_wvalid)
);


wire [IDWID-1:0] merger3_merger4_arid ;
wire [31:0] merger3_merger4_araddr ;
wire [7:0] merger3_merger4_arlen ;
wire [2:0] merger3_merger4_arsize ;
wire [EXTRAS-1:0] merger3_merger4_arextras ;
wire [1:0] merger3_merger4_arburst ;
wire merger3_merger4_arvalid ;
wire merger3_merger4_arready ;
wire [IDWID-1:0] merger3_merger4_rid ;
wire [DWID-1:0] merger3_merger4_rdata ;
wire [1:0] merger3_merger4_rresp ;
wire merger3_merger4_rlast ;
wire merger3_merger4_rvalid ;
wire merger3_merger4_rready ;

wire [IDWID-1:0] merger3_merger4_awid ;
wire [31:0] merger3_merger4_awaddr ;
wire [7:0] merger3_merger4_awlen ;
wire [2:0] merger3_merger4_awsize ;
wire [EXTRAS-1:0] merger3_merger4_awextras ;
wire [1:0] merger3_merger4_awburst ;
wire merger3_merger4_awvalid ;
wire merger3_merger4_awready ;
wire [DWID-1:0] merger3_merger4_wdata ;
wire [WSTRB-1:0] merger3_merger4_wstrb ;
wire merger3_merger4_wlast ;
wire merger3_merger4_wvalid ;
wire merger3_merger4_wready ;
wire [IDWID-1:0] merger3_merger4_bid ;
wire [1:0] merger3_merger4_bresp ;
wire merger3_merger4_bvalid ;
wire merger3_merger4_bready ;


axi_4_merger merger3 (
     .clk(clk),.rst_n(rst_n)
    ,.araddr(merger3_merger4_araddr[31:0])
    ,.arburst(merger3_merger4_arburst[1:0])
    ,.arextras(merger3_merger4_arextras[(EXTRAS - 1):0])
    ,.arid(merger3_merger4_arid)
    ,.arlen(merger3_merger4_arlen)
    ,.arsize(merger3_merger4_arsize)
    ,.arready(merger3_merger4_arready)
    ,.arvalid(merger3_merger4_arvalid)
    ,.awaddr(merger3_merger4_awaddr[31:0])
    ,.awburst(merger3_merger4_awburst[1:0])
    ,.awextras(merger3_merger4_awextras[(EXTRAS - 1):0])
    ,.awid(merger3_merger4_awid)
    ,.awlen(merger3_merger4_awlen)
    ,.awsize(merger3_merger4_awsize)
    ,.awready(merger3_merger4_awready)
    ,.awvalid(merger3_merger4_awvalid)
    ,.bid(merger3_merger4_bid[(IDWID - 1):0])
    ,.bready(merger3_merger4_bready)
    ,.bresp(merger3_merger4_bresp[1:0])
    ,.bvalid(merger3_merger4_bvalid)
    ,.rid(merger3_merger4_rid[(IDWID - 1):0])
    ,.rlast(merger3_merger4_rlast)
    ,.rready(merger3_merger4_rready)
    ,.rresp(merger3_merger4_rresp[1:0])
    ,.rvalid(merger3_merger4_rvalid)
    ,.rdata(merger3_merger4_rdata[(DWID - 1):0])
    ,.wdata(merger3_merger4_wdata[(DWID - 1):0])
    ,.wlast(merger3_merger4_wlast)
    ,.wready(merger3_merger4_wready)
    ,.wstrb(merger3_merger4_wstrb[(WSTRB - 1):0])
    ,.wvalid(merger3_merger4_wvalid)


    ,.a_araddr(mst12_araddr[31:0])
    ,.a_arburst(mst12_arburst[1:0])
    ,.a_arextras(mst12_arextras[(EXTRAS - 1):0])
    ,.a_arid(mst12_arid)
    ,.a_arlen(mst12_arlen)
    ,.a_arsize(mst12_arsize)
    ,.a_arready(mst12_arready)
    ,.a_arvalid(mst12_arvalid)
    ,.a_awaddr(mst12_awaddr[31:0])
    ,.a_awburst(mst12_awburst[1:0])
    ,.a_awextras(mst12_awextras[(EXTRAS - 1):0])
    ,.a_awid(mst12_awid)
    ,.a_awlen(mst12_awlen)
    ,.a_awsize(mst12_awsize)
    ,.a_awready(mst12_awready)
    ,.a_awvalid(mst12_awvalid)
    ,.a_bid(mst12_bid[(IDWID - 1):0])
    ,.a_bready(mst12_bready)
    ,.a_bresp(mst12_bresp[1:0])
    ,.a_bvalid(mst12_bvalid)
    ,.a_rdata(mst12_rdata[(DWID - 1):0])
    ,.a_rid(mst12_rid[(IDWID - 1):0])
    ,.a_rlast(mst12_rlast)
    ,.a_rready(mst12_rready)
    ,.a_rresp(mst12_rresp[1:0])
    ,.a_rvalid(mst12_rvalid)
    ,.a_wdata(mst12_wdata[(DWID - 1):0])
    ,.a_wlast(mst12_wlast)
    ,.a_wready(mst12_wready)
    ,.a_wstrb(mst12_wstrb[(WSTRB - 1):0])
    ,.a_wvalid(mst12_wvalid)

    ,.b_araddr(mst13_araddr[31:0])
    ,.b_arburst(mst13_arburst[1:0])
    ,.b_arextras(mst13_arextras[(EXTRAS - 1):0])
    ,.b_arid(mst13_arid)
    ,.b_arlen(mst13_arlen)
    ,.b_arsize(mst13_arsize)
    ,.b_arready(mst13_arready)
    ,.b_arvalid(mst13_arvalid)
    ,.b_awaddr(mst13_awaddr[31:0])
    ,.b_awburst(mst13_awburst[1:0])
    ,.b_awextras(mst13_awextras[(EXTRAS - 1):0])
    ,.b_awid(mst13_awid)
    ,.b_awlen(mst13_awlen)
    ,.b_awsize(mst13_awsize)
    ,.b_awready(mst13_awready)
    ,.b_awvalid(mst13_awvalid)
    ,.b_bid(mst13_bid[(IDWID - 1):0])
    ,.b_bready(mst13_bready)
    ,.b_bresp(mst13_bresp[1:0])
    ,.b_bvalid(mst13_bvalid)
    ,.b_rdata(mst13_rdata[(DWID - 1):0])
    ,.b_rid(mst13_rid[(IDWID - 1):0])
    ,.b_rlast(mst13_rlast)
    ,.b_rready(mst13_rready)
    ,.b_rresp(mst13_rresp[1:0])
    ,.b_rvalid(mst13_rvalid)
    ,.b_wdata(mst13_wdata[(DWID - 1):0])
    ,.b_wlast(mst13_wlast)
    ,.b_wready(mst13_wready)
    ,.b_wstrb(mst13_wstrb[(WSTRB - 1):0])
    ,.b_wvalid(mst13_wvalid)

    ,.c_araddr(mst14_araddr[31:0])
    ,.c_arburst(mst14_arburst[1:0])
    ,.c_arextras(mst14_arextras[(EXTRAS - 1):0])
    ,.c_arid(mst14_arid)
    ,.c_arlen(mst14_arlen)
    ,.c_arsize(mst14_arsize)
    ,.c_arready(mst14_arready)
    ,.c_arvalid(mst14_arvalid)
    ,.c_awaddr(mst14_awaddr[31:0])
    ,.c_awburst(mst14_awburst[1:0])
    ,.c_awextras(mst14_awextras[(EXTRAS - 1):0])
    ,.c_awid(mst14_awid)
    ,.c_awlen(mst14_awlen)
    ,.c_awsize(mst14_awsize)
    ,.c_awready(mst14_awready)
    ,.c_awvalid(mst14_awvalid)
    ,.c_bid(mst14_bid[(IDWID - 1):0])
    ,.c_bready(mst14_bready)
    ,.c_bresp(mst14_bresp[1:0])
    ,.c_bvalid(mst14_bvalid)
    ,.c_rdata(mst14_rdata[(DWID - 1):0])
    ,.c_rid(mst14_rid[(IDWID - 1):0])
    ,.c_rlast(mst14_rlast)
    ,.c_rready(mst14_rready)
    ,.c_rresp(mst14_rresp[1:0])
    ,.c_rvalid(mst14_rvalid)
    ,.c_wdata(mst14_wdata[(DWID - 1):0])
    ,.c_wlast(mst14_wlast)
    ,.c_wready(mst14_wready)
    ,.c_wstrb(mst14_wstrb[(WSTRB - 1):0])
    ,.c_wvalid(mst14_wvalid)

    ,.d_araddr(mst15_araddr[31:0])
    ,.d_arburst(mst15_arburst[1:0])
    ,.d_arextras(mst15_arextras[(EXTRAS - 1):0])
    ,.d_arid(mst15_arid)
    ,.d_arlen(mst15_arlen)
    ,.d_arsize(mst15_arsize)
    ,.d_arready(mst15_arready)
    ,.d_arvalid(mst15_arvalid)
    ,.d_awaddr(mst15_awaddr[31:0])
    ,.d_awburst(mst15_awburst[1:0])
    ,.d_awextras(mst15_awextras[(EXTRAS - 1):0])
    ,.d_awid(mst15_awid)
    ,.d_awlen(mst15_awlen)
    ,.d_awsize(mst15_awsize)
    ,.d_awready(mst15_awready)
    ,.d_awvalid(mst15_awvalid)
    ,.d_bid(mst15_bid[(IDWID - 1):0])
    ,.d_bready(mst15_bready)
    ,.d_bresp(mst15_bresp[1:0])
    ,.d_bvalid(mst15_bvalid)
    ,.d_rdata(mst15_rdata[(DWID - 1):0])
    ,.d_rid(mst15_rid[(IDWID - 1):0])
    ,.d_rlast(mst15_rlast)
    ,.d_rready(mst15_rready)
    ,.d_rresp(mst15_rresp[1:0])
    ,.d_rvalid(mst15_rvalid)
    ,.d_wdata(mst15_wdata[(DWID - 1):0])
    ,.d_wlast(mst15_wlast)
    ,.d_wready(mst15_wready)
    ,.d_wstrb(mst15_wstrb[(WSTRB - 1):0])
    ,.d_wvalid(mst15_wvalid)
);


wire [IDWID-1:0] merger4_splitter0_arid ;
wire [31:0] merger4_splitter0_araddr ;
wire [7:0] merger4_splitter0_arlen ;
wire [2:0] merger4_splitter0_arsize ;
wire [EXTRAS-1:0] merger4_splitter0_arextras ;
wire [1:0] merger4_splitter0_arburst ;
wire merger4_splitter0_arvalid ;
wire merger4_splitter0_arready ;
wire [IDWID-1:0] merger4_splitter0_rid ;
wire [DWID-1:0] merger4_splitter0_rdata ;
wire [1:0] merger4_splitter0_rresp ;
wire merger4_splitter0_rlast ;
wire merger4_splitter0_rvalid ;
wire merger4_splitter0_rready ;

wire [IDWID-1:0] merger4_splitter0_awid ;
wire [31:0] merger4_splitter0_awaddr ;
wire [7:0] merger4_splitter0_awlen ;
wire [2:0] merger4_splitter0_awsize ;
wire [EXTRAS-1:0] merger4_splitter0_awextras ;
wire [1:0] merger4_splitter0_awburst ;
wire merger4_splitter0_awvalid ;
wire merger4_splitter0_awready ;
wire [DWID-1:0] merger4_splitter0_wdata ;
wire [WSTRB-1:0] merger4_splitter0_wstrb ;
wire merger4_splitter0_wlast ;
wire merger4_splitter0_wvalid ;
wire merger4_splitter0_wready ;
wire [IDWID-1:0] merger4_splitter0_bid ;
wire [1:0] merger4_splitter0_bresp ;
wire merger4_splitter0_bvalid ;
wire merger4_splitter0_bready ;


axi_4_merger merger4 (
     .clk(clk),.rst_n(rst_n)
    ,.araddr(merger4_splitter0_araddr[31:0])
    ,.arburst(merger4_splitter0_arburst[1:0])
    ,.arextras(merger4_splitter0_arextras[(EXTRAS - 1):0])
    ,.arid(merger4_splitter0_arid)
    ,.arlen(merger4_splitter0_arlen)
    ,.arsize(merger4_splitter0_arsize)
    ,.arready(merger4_splitter0_arready)
    ,.arvalid(merger4_splitter0_arvalid)
    ,.awaddr(merger4_splitter0_awaddr[31:0])
    ,.awburst(merger4_splitter0_awburst[1:0])
    ,.awextras(merger4_splitter0_awextras[(EXTRAS - 1):0])
    ,.awid(merger4_splitter0_awid)
    ,.awlen(merger4_splitter0_awlen)
    ,.awsize(merger4_splitter0_awsize)
    ,.awready(merger4_splitter0_awready)
    ,.awvalid(merger4_splitter0_awvalid)
    ,.bid(merger4_splitter0_bid[(IDWID - 1):0])
    ,.bready(merger4_splitter0_bready)
    ,.bresp(merger4_splitter0_bresp[1:0])
    ,.bvalid(merger4_splitter0_bvalid)
    ,.rid(merger4_splitter0_rid[(IDWID - 1):0])
    ,.rlast(merger4_splitter0_rlast)
    ,.rready(merger4_splitter0_rready)
    ,.rresp(merger4_splitter0_rresp[1:0])
    ,.rvalid(merger4_splitter0_rvalid)
    ,.rdata(merger4_splitter0_rdata[(DWID - 1):0])
    ,.wdata(merger4_splitter0_wdata[(DWID - 1):0])
    ,.wlast(merger4_splitter0_wlast)
    ,.wready(merger4_splitter0_wready)
    ,.wstrb(merger4_splitter0_wstrb[(WSTRB - 1):0])
    ,.wvalid(merger4_splitter0_wvalid)


    ,.a_araddr(merger0_merger4_araddr[31:0])
    ,.a_arburst(merger0_merger4_arburst[1:0])
    ,.a_arextras(merger0_merger4_arextras[(EXTRAS - 1):0])
    ,.a_arid(merger0_merger4_arid)
    ,.a_arlen(merger0_merger4_arlen)
    ,.a_arsize(merger0_merger4_arsize)
    ,.a_arready(merger0_merger4_arready)
    ,.a_arvalid(merger0_merger4_arvalid)
    ,.a_awaddr(merger0_merger4_awaddr[31:0])
    ,.a_awburst(merger0_merger4_awburst[1:0])
    ,.a_awextras(merger0_merger4_awextras[(EXTRAS - 1):0])
    ,.a_awid(merger0_merger4_awid)
    ,.a_awlen(merger0_merger4_awlen)
    ,.a_awsize(merger0_merger4_awsize)
    ,.a_awready(merger0_merger4_awready)
    ,.a_awvalid(merger0_merger4_awvalid)
    ,.a_bid(merger0_merger4_bid[(IDWID - 1):0])
    ,.a_bready(merger0_merger4_bready)
    ,.a_bresp(merger0_merger4_bresp[1:0])
    ,.a_bvalid(merger0_merger4_bvalid)
    ,.a_rdata(merger0_merger4_rdata[(DWID - 1):0])
    ,.a_rid(merger0_merger4_rid[(IDWID - 1):0])
    ,.a_rlast(merger0_merger4_rlast)
    ,.a_rready(merger0_merger4_rready)
    ,.a_rresp(merger0_merger4_rresp[1:0])
    ,.a_rvalid(merger0_merger4_rvalid)
    ,.a_wdata(merger0_merger4_wdata[(DWID - 1):0])
    ,.a_wlast(merger0_merger4_wlast)
    ,.a_wready(merger0_merger4_wready)
    ,.a_wstrb(merger0_merger4_wstrb[(WSTRB - 1):0])
    ,.a_wvalid(merger0_merger4_wvalid)

    ,.b_araddr(merger1_merger4_araddr[31:0])
    ,.b_arburst(merger1_merger4_arburst[1:0])
    ,.b_arextras(merger1_merger4_arextras[(EXTRAS - 1):0])
    ,.b_arid(merger1_merger4_arid)
    ,.b_arlen(merger1_merger4_arlen)
    ,.b_arsize(merger1_merger4_arsize)
    ,.b_arready(merger1_merger4_arready)
    ,.b_arvalid(merger1_merger4_arvalid)
    ,.b_awaddr(merger1_merger4_awaddr[31:0])
    ,.b_awburst(merger1_merger4_awburst[1:0])
    ,.b_awextras(merger1_merger4_awextras[(EXTRAS - 1):0])
    ,.b_awid(merger1_merger4_awid)
    ,.b_awlen(merger1_merger4_awlen)
    ,.b_awsize(merger1_merger4_awsize)
    ,.b_awready(merger1_merger4_awready)
    ,.b_awvalid(merger1_merger4_awvalid)
    ,.b_bid(merger1_merger4_bid[(IDWID - 1):0])
    ,.b_bready(merger1_merger4_bready)
    ,.b_bresp(merger1_merger4_bresp[1:0])
    ,.b_bvalid(merger1_merger4_bvalid)
    ,.b_rdata(merger1_merger4_rdata[(DWID - 1):0])
    ,.b_rid(merger1_merger4_rid[(IDWID - 1):0])
    ,.b_rlast(merger1_merger4_rlast)
    ,.b_rready(merger1_merger4_rready)
    ,.b_rresp(merger1_merger4_rresp[1:0])
    ,.b_rvalid(merger1_merger4_rvalid)
    ,.b_wdata(merger1_merger4_wdata[(DWID - 1):0])
    ,.b_wlast(merger1_merger4_wlast)
    ,.b_wready(merger1_merger4_wready)
    ,.b_wstrb(merger1_merger4_wstrb[(WSTRB - 1):0])
    ,.b_wvalid(merger1_merger4_wvalid)

    ,.c_araddr(merger2_merger4_araddr[31:0])
    ,.c_arburst(merger2_merger4_arburst[1:0])
    ,.c_arextras(merger2_merger4_arextras[(EXTRAS - 1):0])
    ,.c_arid(merger2_merger4_arid)
    ,.c_arlen(merger2_merger4_arlen)
    ,.c_arsize(merger2_merger4_arsize)
    ,.c_arready(merger2_merger4_arready)
    ,.c_arvalid(merger2_merger4_arvalid)
    ,.c_awaddr(merger2_merger4_awaddr[31:0])
    ,.c_awburst(merger2_merger4_awburst[1:0])
    ,.c_awextras(merger2_merger4_awextras[(EXTRAS - 1):0])
    ,.c_awid(merger2_merger4_awid)
    ,.c_awlen(merger2_merger4_awlen)
    ,.c_awsize(merger2_merger4_awsize)
    ,.c_awready(merger2_merger4_awready)
    ,.c_awvalid(merger2_merger4_awvalid)
    ,.c_bid(merger2_merger4_bid[(IDWID - 1):0])
    ,.c_bready(merger2_merger4_bready)
    ,.c_bresp(merger2_merger4_bresp[1:0])
    ,.c_bvalid(merger2_merger4_bvalid)
    ,.c_rdata(merger2_merger4_rdata[(DWID - 1):0])
    ,.c_rid(merger2_merger4_rid[(IDWID - 1):0])
    ,.c_rlast(merger2_merger4_rlast)
    ,.c_rready(merger2_merger4_rready)
    ,.c_rresp(merger2_merger4_rresp[1:0])
    ,.c_rvalid(merger2_merger4_rvalid)
    ,.c_wdata(merger2_merger4_wdata[(DWID - 1):0])
    ,.c_wlast(merger2_merger4_wlast)
    ,.c_wready(merger2_merger4_wready)
    ,.c_wstrb(merger2_merger4_wstrb[(WSTRB - 1):0])
    ,.c_wvalid(merger2_merger4_wvalid)

    ,.d_araddr(merger3_merger4_araddr[31:0])
    ,.d_arburst(merger3_merger4_arburst[1:0])
    ,.d_arextras(merger3_merger4_arextras[(EXTRAS - 1):0])
    ,.d_arid(merger3_merger4_arid)
    ,.d_arlen(merger3_merger4_arlen)
    ,.d_arsize(merger3_merger4_arsize)
    ,.d_arready(merger3_merger4_arready)
    ,.d_arvalid(merger3_merger4_arvalid)
    ,.d_awaddr(merger3_merger4_awaddr[31:0])
    ,.d_awburst(merger3_merger4_awburst[1:0])
    ,.d_awextras(merger3_merger4_awextras[(EXTRAS - 1):0])
    ,.d_awid(merger3_merger4_awid)
    ,.d_awlen(merger3_merger4_awlen)
    ,.d_awsize(merger3_merger4_awsize)
    ,.d_awready(merger3_merger4_awready)
    ,.d_awvalid(merger3_merger4_awvalid)
    ,.d_bid(merger3_merger4_bid[(IDWID - 1):0])
    ,.d_bready(merger3_merger4_bready)
    ,.d_bresp(merger3_merger4_bresp[1:0])
    ,.d_bvalid(merger3_merger4_bvalid)
    ,.d_rdata(merger3_merger4_rdata[(DWID - 1):0])
    ,.d_rid(merger3_merger4_rid[(IDWID - 1):0])
    ,.d_rlast(merger3_merger4_rlast)
    ,.d_rready(merger3_merger4_rready)
    ,.d_rresp(merger3_merger4_rresp[1:0])
    ,.d_rvalid(merger3_merger4_rvalid)
    ,.d_wdata(merger3_merger4_wdata[(DWID - 1):0])
    ,.d_wlast(merger3_merger4_wlast)
    ,.d_wready(merger3_merger4_wready)
    ,.d_wstrb(merger3_merger4_wstrb[(WSTRB - 1):0])
    ,.d_wvalid(merger3_merger4_wvalid)
);


axi_4_splitter splitter0 (
     .clk(clk) ,.rst_n(rst_n)

    ,.araddr(merger4_splitter0_araddr[31:0])
    ,.arburst(merger4_splitter0_arburst[1:0])
    ,.arextras(merger4_splitter0_arextras[(EXTRAS - 1):0])
    ,.arid(merger4_splitter0_arid)
    ,.arlen(merger4_splitter0_arlen)
    ,.arsize(merger4_splitter0_arsize)
    ,.arready(merger4_splitter0_arready)
    ,.arvalid(merger4_splitter0_arvalid)
    ,.awaddr(merger4_splitter0_awaddr[31:0])
    ,.awburst(merger4_splitter0_awburst[1:0])
    ,.awextras(merger4_splitter0_awextras[(EXTRAS - 1):0])
    ,.awid(merger4_splitter0_awid)
    ,.awlen(merger4_splitter0_awlen)
    ,.awsize(merger4_splitter0_awsize)
    ,.awready(merger4_splitter0_awready)
    ,.awvalid(merger4_splitter0_awvalid)
    ,.bid(merger4_splitter0_bid[(IDWID - 1):0])
    ,.bready(merger4_splitter0_bready)
    ,.bresp(merger4_splitter0_bresp[1:0])
    ,.bvalid(merger4_splitter0_bvalid)
    ,.rdata(merger4_splitter0_rdata[(DWID - 1):0])
    ,.rid(merger4_splitter0_rid[(IDWID - 1):0])
    ,.rlast(merger4_splitter0_rlast)
    ,.rready(merger4_splitter0_rready)
    ,.rresp(merger4_splitter0_rresp[1:0])
    ,.rvalid(merger4_splitter0_rvalid)
    ,.wdata(merger4_splitter0_wdata[(DWID - 1):0])
    ,.wlast(merger4_splitter0_wlast)
    ,.wready(merger4_splitter0_wready)
    ,.wstrb(merger4_splitter0_wstrb[(WSTRB - 1):0])
    ,.wvalid(merger4_splitter0_wvalid)

    ,.a_araddr(slv0_araddr[31:0])
    ,.a_arburst(slv0_arburst[1:0])
    ,.a_arextras(slv0_arextras[(EXTRAS - 1):0])
    ,.a_arid(slv0_arid)
    ,.a_arlen(slv0_arlen)
    ,.a_arsize(slv0_arsize)
    ,.a_arready(slv0_arready)
    ,.a_arvalid(slv0_arvalid)
    ,.a_awaddr(slv0_awaddr[31:0])
    ,.a_awburst(slv0_awburst[1:0])
    ,.a_awextras(slv0_awextras[(EXTRAS - 1):0])
    ,.a_awid(slv0_awid)
    ,.a_awlen(slv0_awlen)
    ,.a_awsize(slv0_awsize)
    ,.a_awready(slv0_awready)
    ,.a_awvalid(slv0_awvalid)
    ,.a_bid(slv0_bid[(IDWID - 1):0])
    ,.a_bready(slv0_bready)
    ,.a_bresp(slv0_bresp[1:0])
    ,.a_bvalid(slv0_bvalid)
    ,.a_rdata(slv0_rdata[(DWID - 1):0])
    ,.a_rid(slv0_rid[(IDWID - 1):0])
    ,.a_rlast(slv0_rlast)
    ,.a_rready(slv0_rready)
    ,.a_rresp(slv0_rresp[1:0])
    ,.a_rvalid(slv0_rvalid)
    ,.a_wdata(slv0_wdata[(DWID - 1):0])
    ,.a_wlast(slv0_wlast)
    ,.a_wready(slv0_wready)
    ,.a_wstrb(slv0_wstrb[(WSTRB - 1):0])
    ,.a_wvalid(slv0_wvalid)
    ,.b_araddr(slv1_araddr[31:0])
    ,.b_arburst(slv1_arburst[1:0])
    ,.b_arextras(slv1_arextras[(EXTRAS - 1):0])
    ,.b_arid(slv1_arid)
    ,.b_arlen(slv1_arlen)
    ,.b_arsize(slv1_arsize)
    ,.b_arready(slv1_arready)
    ,.b_arvalid(slv1_arvalid)
    ,.b_awaddr(slv1_awaddr[31:0])
    ,.b_awburst(slv1_awburst[1:0])
    ,.b_awextras(slv1_awextras[(EXTRAS - 1):0])
    ,.b_awid(slv1_awid)
    ,.b_awlen(slv1_awlen)
    ,.b_awsize(slv1_awsize)
    ,.b_awready(slv1_awready)
    ,.b_awvalid(slv1_awvalid)
    ,.b_bid(slv1_bid[(IDWID - 1):0])
    ,.b_bready(slv1_bready)
    ,.b_bresp(slv1_bresp[1:0])
    ,.b_bvalid(slv1_bvalid)
    ,.b_rdata(slv1_rdata[(DWID - 1):0])
    ,.b_rid(slv1_rid[(IDWID - 1):0])
    ,.b_rlast(slv1_rlast)
    ,.b_rready(slv1_rready)
    ,.b_rresp(slv1_rresp[1:0])
    ,.b_rvalid(slv1_rvalid)
    ,.b_wdata(slv1_wdata[(DWID - 1):0])
    ,.b_wlast(slv1_wlast)
    ,.b_wready(slv1_wready)
    ,.b_wstrb(slv1_wstrb[(WSTRB - 1):0])
    ,.b_wvalid(slv1_wvalid)
    ,.c_araddr(slv2_araddr[31:0])
    ,.c_arburst(slv2_arburst[1:0])
    ,.c_arextras(slv2_arextras[(EXTRAS - 1):0])
    ,.c_arid(slv2_arid)
    ,.c_arlen(slv2_arlen)
    ,.c_arsize(slv2_arsize)
    ,.c_arready(slv2_arready)
    ,.c_arvalid(slv2_arvalid)
    ,.c_awaddr(slv2_awaddr[31:0])
    ,.c_awburst(slv2_awburst[1:0])
    ,.c_awextras(slv2_awextras[(EXTRAS - 1):0])
    ,.c_awid(slv2_awid)
    ,.c_awlen(slv2_awlen)
    ,.c_awsize(slv2_awsize)
    ,.c_awready(slv2_awready)
    ,.c_awvalid(slv2_awvalid)
    ,.c_bid(slv2_bid[(IDWID - 1):0])
    ,.c_bready(slv2_bready)
    ,.c_bresp(slv2_bresp[1:0])
    ,.c_bvalid(slv2_bvalid)
    ,.c_rdata(slv2_rdata[(DWID - 1):0])
    ,.c_rid(slv2_rid[(IDWID - 1):0])
    ,.c_rlast(slv2_rlast)
    ,.c_rready(slv2_rready)
    ,.c_rresp(slv2_rresp[1:0])
    ,.c_rvalid(slv2_rvalid)
    ,.c_wdata(slv2_wdata[(DWID - 1):0])
    ,.c_wlast(slv2_wlast)
    ,.c_wready(slv2_wready)
    ,.c_wstrb(slv2_wstrb[(WSTRB - 1):0])
    ,.c_wvalid(slv2_wvalid)
    ,.d_araddr(slv3_araddr[31:0])
    ,.d_arburst(slv3_arburst[1:0])
    ,.d_arextras(slv3_arextras[(EXTRAS - 1):0])
    ,.d_arid(slv3_arid[(IDWID - 1):0])
    ,.d_arlen(slv3_arlen[7:0])
    ,.d_arsize(slv3_arsize)
    ,.d_arready(slv3_arready)
    ,.d_arvalid(slv3_arvalid)
    ,.d_awaddr(slv3_awaddr[31:0])
    ,.d_awburst(slv3_awburst[1:0])
    ,.d_awextras(slv3_awextras[(EXTRAS - 1):0])
    ,.d_awid(slv3_awid)
    ,.d_awlen(slv3_awlen)
    ,.d_awsize(slv3_awsize)
    ,.d_awready(slv3_awready)
    ,.d_awvalid(slv3_awvalid)
    ,.d_bid(slv3_bid[(IDWID - 1):0])
    ,.d_bready(slv3_bready)
    ,.d_bresp(slv3_bresp[1:0])
    ,.d_bvalid(slv3_bvalid)
    ,.d_rdata(slv3_rdata[(DWID - 1):0])
    ,.d_rid(slv3_rid[(IDWID - 1):0])
    ,.d_rlast(slv3_rlast)
    ,.d_rready(slv3_rready)
    ,.d_rresp(slv3_rresp[1:0])
    ,.d_rvalid(slv3_rvalid)
    ,.d_wdata(slv3_wdata[(DWID - 1):0])
    ,.d_wlast(slv3_wlast)
    ,.d_wready(slv3_wready)
    ,.d_wstrb(slv3_wstrb[(WSTRB - 1):0])
    ,.d_wvalid(slv3_wvalid)

);
endmodule
