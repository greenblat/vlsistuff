module sintab(input [10:0] addr,output reg [15:0] out);
always @* begin
    case (addr)
        0 : out = 0;
        1 : out = 100;
        2 : out = 201;
        3 : out = 301;
        4 : out = 402;
        5 : out = 502;
        6 : out = 603;
        7 : out = 703;
        8 : out = 804;
        9 : out = 904;
        10 : out = 1005;
        11 : out = 1105;
        12 : out = 1206;
        13 : out = 1306;
        14 : out = 1406;
        15 : out = 1507;
        16 : out = 1607;
        17 : out = 1708;
        18 : out = 1808;
        19 : out = 1908;
        20 : out = 2009;
        21 : out = 2109;
        22 : out = 2209;
        23 : out = 2310;
        24 : out = 2410;
        25 : out = 2510;
        26 : out = 2610;
        27 : out = 2711;
        28 : out = 2811;
        29 : out = 2911;
        30 : out = 3011;
        31 : out = 3111;
        32 : out = 3211;
        33 : out = 3311;
        34 : out = 3411;
        35 : out = 3511;
        36 : out = 3611;
        37 : out = 3711;
        38 : out = 3811;
        39 : out = 3911;
        40 : out = 4011;
        41 : out = 4110;
        42 : out = 4210;
        43 : out = 4310;
        44 : out = 4409;
        45 : out = 4509;
        46 : out = 4608;
        47 : out = 4708;
        48 : out = 4807;
        49 : out = 4907;
        50 : out = 5006;
        51 : out = 5106;
        52 : out = 5205;
        53 : out = 5304;
        54 : out = 5403;
        55 : out = 5502;
        56 : out = 5601;
        57 : out = 5700;
        58 : out = 5799;
        59 : out = 5898;
        60 : out = 5997;
        61 : out = 6096;
        62 : out = 6195;
        63 : out = 6293;
        64 : out = 6392;
        65 : out = 6491;
        66 : out = 6589;
        67 : out = 6688;
        68 : out = 6786;
        69 : out = 6884;
        70 : out = 6982;
        71 : out = 7081;
        72 : out = 7179;
        73 : out = 7277;
        74 : out = 7375;
        75 : out = 7473;
        76 : out = 7571;
        77 : out = 7668;
        78 : out = 7766;
        79 : out = 7864;
        80 : out = 7961;
        81 : out = 8059;
        82 : out = 8156;
        83 : out = 8253;
        84 : out = 8351;
        85 : out = 8448;
        86 : out = 8545;
        87 : out = 8642;
        88 : out = 8739;
        89 : out = 8836;
        90 : out = 8932;
        91 : out = 9029;
        92 : out = 9126;
        93 : out = 9222;
        94 : out = 9319;
        95 : out = 9415;
        96 : out = 9511;
        97 : out = 9607;
        98 : out = 9703;
        99 : out = 9799;
        100 : out = 9895;
        101 : out = 9991;
        102 : out = 10087;
        103 : out = 10182;
        104 : out = 10278;
        105 : out = 10373;
        106 : out = 10469;
        107 : out = 10564;
        108 : out = 10659;
        109 : out = 10754;
        110 : out = 10849;
        111 : out = 10944;
        112 : out = 11038;
        113 : out = 11133;
        114 : out = 11227;
        115 : out = 11322;
        116 : out = 11416;
        117 : out = 11510;
        118 : out = 11604;
        119 : out = 11698;
        120 : out = 11792;
        121 : out = 11886;
        122 : out = 11980;
        123 : out = 12073;
        124 : out = 12166;
        125 : out = 12260;
        126 : out = 12353;
        127 : out = 12446;
        128 : out = 12539;
        129 : out = 12632;
        130 : out = 12724;
        131 : out = 12817;
        132 : out = 12909;
        133 : out = 13002;
        134 : out = 13094;
        135 : out = 13186;
        136 : out = 13278;
        137 : out = 13370;
        138 : out = 13462;
        139 : out = 13553;
        140 : out = 13645;
        141 : out = 13736;
        142 : out = 13827;
        143 : out = 13918;
        144 : out = 14009;
        145 : out = 14100;
        146 : out = 14191;
        147 : out = 14281;
        148 : out = 14372;
        149 : out = 14462;
        150 : out = 14552;
        151 : out = 14642;
        152 : out = 14732;
        153 : out = 14822;
        154 : out = 14911;
        155 : out = 15001;
        156 : out = 15090;
        157 : out = 15179;
        158 : out = 15268;
        159 : out = 15357;
        160 : out = 15446;
        161 : out = 15534;
        162 : out = 15623;
        163 : out = 15711;
        164 : out = 15799;
        165 : out = 15887;
        166 : out = 15975;
        167 : out = 16063;
        168 : out = 16150;
        169 : out = 16238;
        170 : out = 16325;
        171 : out = 16412;
        172 : out = 16499;
        173 : out = 16586;
        174 : out = 16672;
        175 : out = 16759;
        176 : out = 16845;
        177 : out = 16931;
        178 : out = 17017;
        179 : out = 17103;
        180 : out = 17189;
        181 : out = 17274;
        182 : out = 17360;
        183 : out = 17445;
        184 : out = 17530;
        185 : out = 17615;
        186 : out = 17699;
        187 : out = 17784;
        188 : out = 17868;
        189 : out = 17952;
        190 : out = 18036;
        191 : out = 18120;
        192 : out = 18204;
        193 : out = 18287;
        194 : out = 18371;
        195 : out = 18454;
        196 : out = 18537;
        197 : out = 18620;
        198 : out = 18702;
        199 : out = 18785;
        200 : out = 18867;
        201 : out = 18949;
        202 : out = 19031;
        203 : out = 19113;
        204 : out = 19194;
        205 : out = 19276;
        206 : out = 19357;
        207 : out = 19438;
        208 : out = 19519;
        209 : out = 19599;
        210 : out = 19680;
        211 : out = 19760;
        212 : out = 19840;
        213 : out = 19920;
        214 : out = 20000;
        215 : out = 20079;
        216 : out = 20159;
        217 : out = 20238;
        218 : out = 20317;
        219 : out = 20396;
        220 : out = 20474;
        221 : out = 20553;
        222 : out = 20631;
        223 : out = 20709;
        224 : out = 20787;
        225 : out = 20864;
        226 : out = 20942;
        227 : out = 21019;
        228 : out = 21096;
        229 : out = 21173;
        230 : out = 21249;
        231 : out = 21326;
        232 : out = 21402;
        233 : out = 21478;
        234 : out = 21554;
        235 : out = 21629;
        236 : out = 21705;
        237 : out = 21780;
        238 : out = 21855;
        239 : out = 21930;
        240 : out = 22004;
        241 : out = 22079;
        242 : out = 22153;
        243 : out = 22227;
        244 : out = 22301;
        245 : out = 22374;
        246 : out = 22448;
        247 : out = 22521;
        248 : out = 22594;
        249 : out = 22666;
        250 : out = 22739;
        251 : out = 22811;
        252 : out = 22883;
        253 : out = 22955;
        254 : out = 23027;
        255 : out = 23098;
        256 : out = 23169;
        257 : out = 23240;
        258 : out = 23311;
        259 : out = 23382;
        260 : out = 23452;
        261 : out = 23522;
        262 : out = 23592;
        263 : out = 23661;
        264 : out = 23731;
        265 : out = 23800;
        266 : out = 23869;
        267 : out = 23938;
        268 : out = 24006;
        269 : out = 24075;
        270 : out = 24143;
        271 : out = 24211;
        272 : out = 24278;
        273 : out = 24346;
        274 : out = 24413;
        275 : out = 24480;
        276 : out = 24546;
        277 : out = 24613;
        278 : out = 24679;
        279 : out = 24745;
        280 : out = 24811;
        281 : out = 24877;
        282 : out = 24942;
        283 : out = 25007;
        284 : out = 25072;
        285 : out = 25136;
        286 : out = 25201;
        287 : out = 25265;
        288 : out = 25329;
        289 : out = 25392;
        290 : out = 25456;
        291 : out = 25519;
        292 : out = 25582;
        293 : out = 25645;
        294 : out = 25707;
        295 : out = 25769;
        296 : out = 25831;
        297 : out = 25893;
        298 : out = 25954;
        299 : out = 26016;
        300 : out = 26077;
        301 : out = 26137;
        302 : out = 26198;
        303 : out = 26258;
        304 : out = 26318;
        305 : out = 26378;
        306 : out = 26437;
        307 : out = 26497;
        308 : out = 26556;
        309 : out = 26615;
        310 : out = 26673;
        311 : out = 26731;
        312 : out = 26789;
        313 : out = 26847;
        314 : out = 26905;
        315 : out = 26962;
        316 : out = 27019;
        317 : out = 27076;
        318 : out = 27132;
        319 : out = 27188;
        320 : out = 27244;
        321 : out = 27300;
        322 : out = 27355;
        323 : out = 27411;
        324 : out = 27466;
        325 : out = 27520;
        326 : out = 27575;
        327 : out = 27629;
        328 : out = 27683;
        329 : out = 27736;
        330 : out = 27790;
        331 : out = 27843;
        332 : out = 27896;
        333 : out = 27948;
        334 : out = 28001;
        335 : out = 28053;
        336 : out = 28105;
        337 : out = 28156;
        338 : out = 28208;
        339 : out = 28259;
        340 : out = 28309;
        341 : out = 28360;
        342 : out = 28410;
        343 : out = 28460;
        344 : out = 28510;
        345 : out = 28559;
        346 : out = 28608;
        347 : out = 28657;
        348 : out = 28706;
        349 : out = 28754;
        350 : out = 28802;
        351 : out = 28850;
        352 : out = 28897;
        353 : out = 28945;
        354 : out = 28992;
        355 : out = 29038;
        356 : out = 29085;
        357 : out = 29131;
        358 : out = 29177;
        359 : out = 29222;
        360 : out = 29268;
        361 : out = 29313;
        362 : out = 29358;
        363 : out = 29402;
        364 : out = 29446;
        365 : out = 29490;
        366 : out = 29534;
        367 : out = 29577;
        368 : out = 29621;
        369 : out = 29663;
        370 : out = 29706;
        371 : out = 29748;
        372 : out = 29790;
        373 : out = 29832;
        374 : out = 29873;
        375 : out = 29915;
        376 : out = 29955;
        377 : out = 29996;
        378 : out = 30036;
        379 : out = 30076;
        380 : out = 30116;
        381 : out = 30156;
        382 : out = 30195;
        383 : out = 30234;
        384 : out = 30272;
        385 : out = 30311;
        386 : out = 30349;
        387 : out = 30386;
        388 : out = 30424;
        389 : out = 30461;
        390 : out = 30498;
        391 : out = 30535;
        392 : out = 30571;
        393 : out = 30607;
        394 : out = 30643;
        395 : out = 30678;
        396 : out = 30713;
        397 : out = 30748;
        398 : out = 30783;
        399 : out = 30817;
        400 : out = 30851;
        401 : out = 30885;
        402 : out = 30918;
        403 : out = 30951;
        404 : out = 30984;
        405 : out = 31017;
        406 : out = 31049;
        407 : out = 31081;
        408 : out = 31113;
        409 : out = 31144;
        410 : out = 31175;
        411 : out = 31206;
        412 : out = 31236;
        413 : out = 31267;
        414 : out = 31297;
        415 : out = 31326;
        416 : out = 31356;
        417 : out = 31385;
        418 : out = 31413;
        419 : out = 31442;
        420 : out = 31470;
        421 : out = 31498;
        422 : out = 31525;
        423 : out = 31553;
        424 : out = 31580;
        425 : out = 31606;
        426 : out = 31633;
        427 : out = 31659;
        428 : out = 31684;
        429 : out = 31710;
        430 : out = 31735;
        431 : out = 31760;
        432 : out = 31785;
        433 : out = 31809;
        434 : out = 31833;
        435 : out = 31856;
        436 : out = 31880;
        437 : out = 31903;
        438 : out = 31926;
        439 : out = 31948;
        440 : out = 31970;
        441 : out = 31992;
        442 : out = 32014;
        443 : out = 32035;
        444 : out = 32056;
        445 : out = 32077;
        446 : out = 32097;
        447 : out = 32117;
        448 : out = 32137;
        449 : out = 32156;
        450 : out = 32176;
        451 : out = 32194;
        452 : out = 32213;
        453 : out = 32231;
        454 : out = 32249;
        455 : out = 32267;
        456 : out = 32284;
        457 : out = 32301;
        458 : out = 32318;
        459 : out = 32334;
        460 : out = 32350;
        461 : out = 32366;
        462 : out = 32382;
        463 : out = 32397;
        464 : out = 32412;
        465 : out = 32426;
        466 : out = 32441;
        467 : out = 32455;
        468 : out = 32468;
        469 : out = 32482;
        470 : out = 32495;
        471 : out = 32508;
        472 : out = 32520;
        473 : out = 32532;
        474 : out = 32544;
        475 : out = 32556;
        476 : out = 32567;
        477 : out = 32578;
        478 : out = 32588;
        479 : out = 32599;
        480 : out = 32609;
        481 : out = 32618;
        482 : out = 32628;
        483 : out = 32637;
        484 : out = 32646;
        485 : out = 32654;
        486 : out = 32662;
        487 : out = 32670;
        488 : out = 32678;
        489 : out = 32685;
        490 : out = 32692;
        491 : out = 32699;
        492 : out = 32705;
        493 : out = 32711;
        494 : out = 32717;
        495 : out = 32722;
        496 : out = 32727;
        497 : out = 32732;
        498 : out = 32736;
        499 : out = 32740;
        500 : out = 32744;
        501 : out = 32748;
        502 : out = 32751;
        503 : out = 32754;
        504 : out = 32757;
        505 : out = 32759;
        506 : out = 32761;
        507 : out = 32763;
        508 : out = 32764;
        509 : out = 32765;
        510 : out = 32766;
        511 : out = 32766;
        512 : out = 32767;
        513 : out = 32766;
        514 : out = 32766;
        515 : out = 32765;
        516 : out = 32764;
        517 : out = 32763;
        518 : out = 32761;
        519 : out = 32759;
        520 : out = 32757;
        521 : out = 32754;
        522 : out = 32751;
        523 : out = 32748;
        524 : out = 32744;
        525 : out = 32740;
        526 : out = 32736;
        527 : out = 32732;
        528 : out = 32727;
        529 : out = 32722;
        530 : out = 32717;
        531 : out = 32711;
        532 : out = 32705;
        533 : out = 32699;
        534 : out = 32692;
        535 : out = 32685;
        536 : out = 32678;
        537 : out = 32670;
        538 : out = 32662;
        539 : out = 32654;
        540 : out = 32646;
        541 : out = 32637;
        542 : out = 32628;
        543 : out = 32618;
        544 : out = 32609;
        545 : out = 32599;
        546 : out = 32588;
        547 : out = 32578;
        548 : out = 32567;
        549 : out = 32556;
        550 : out = 32544;
        551 : out = 32532;
        552 : out = 32520;
        553 : out = 32508;
        554 : out = 32495;
        555 : out = 32482;
        556 : out = 32468;
        557 : out = 32455;
        558 : out = 32441;
        559 : out = 32426;
        560 : out = 32412;
        561 : out = 32397;
        562 : out = 32382;
        563 : out = 32366;
        564 : out = 32350;
        565 : out = 32334;
        566 : out = 32318;
        567 : out = 32301;
        568 : out = 32284;
        569 : out = 32267;
        570 : out = 32249;
        571 : out = 32231;
        572 : out = 32213;
        573 : out = 32194;
        574 : out = 32176;
        575 : out = 32156;
        576 : out = 32137;
        577 : out = 32117;
        578 : out = 32097;
        579 : out = 32077;
        580 : out = 32056;
        581 : out = 32035;
        582 : out = 32014;
        583 : out = 31992;
        584 : out = 31970;
        585 : out = 31948;
        586 : out = 31926;
        587 : out = 31903;
        588 : out = 31880;
        589 : out = 31856;
        590 : out = 31833;
        591 : out = 31809;
        592 : out = 31785;
        593 : out = 31760;
        594 : out = 31735;
        595 : out = 31710;
        596 : out = 31684;
        597 : out = 31659;
        598 : out = 31633;
        599 : out = 31606;
        600 : out = 31580;
        601 : out = 31553;
        602 : out = 31525;
        603 : out = 31498;
        604 : out = 31470;
        605 : out = 31442;
        606 : out = 31413;
        607 : out = 31385;
        608 : out = 31356;
        609 : out = 31326;
        610 : out = 31297;
        611 : out = 31267;
        612 : out = 31236;
        613 : out = 31206;
        614 : out = 31175;
        615 : out = 31144;
        616 : out = 31113;
        617 : out = 31081;
        618 : out = 31049;
        619 : out = 31017;
        620 : out = 30984;
        621 : out = 30951;
        622 : out = 30918;
        623 : out = 30885;
        624 : out = 30851;
        625 : out = 30817;
        626 : out = 30783;
        627 : out = 30748;
        628 : out = 30713;
        629 : out = 30678;
        630 : out = 30643;
        631 : out = 30607;
        632 : out = 30571;
        633 : out = 30535;
        634 : out = 30498;
        635 : out = 30461;
        636 : out = 30424;
        637 : out = 30386;
        638 : out = 30349;
        639 : out = 30311;
        640 : out = 30272;
        641 : out = 30234;
        642 : out = 30195;
        643 : out = 30156;
        644 : out = 30116;
        645 : out = 30076;
        646 : out = 30036;
        647 : out = 29996;
        648 : out = 29955;
        649 : out = 29915;
        650 : out = 29873;
        651 : out = 29832;
        652 : out = 29790;
        653 : out = 29748;
        654 : out = 29706;
        655 : out = 29663;
        656 : out = 29621;
        657 : out = 29577;
        658 : out = 29534;
        659 : out = 29490;
        660 : out = 29446;
        661 : out = 29402;
        662 : out = 29358;
        663 : out = 29313;
        664 : out = 29268;
        665 : out = 29222;
        666 : out = 29177;
        667 : out = 29131;
        668 : out = 29085;
        669 : out = 29038;
        670 : out = 28992;
        671 : out = 28945;
        672 : out = 28897;
        673 : out = 28850;
        674 : out = 28802;
        675 : out = 28754;
        676 : out = 28706;
        677 : out = 28657;
        678 : out = 28608;
        679 : out = 28559;
        680 : out = 28510;
        681 : out = 28460;
        682 : out = 28410;
        683 : out = 28360;
        684 : out = 28309;
        685 : out = 28259;
        686 : out = 28208;
        687 : out = 28156;
        688 : out = 28105;
        689 : out = 28053;
        690 : out = 28001;
        691 : out = 27948;
        692 : out = 27896;
        693 : out = 27843;
        694 : out = 27790;
        695 : out = 27736;
        696 : out = 27683;
        697 : out = 27629;
        698 : out = 27575;
        699 : out = 27520;
        700 : out = 27466;
        701 : out = 27411;
        702 : out = 27355;
        703 : out = 27300;
        704 : out = 27244;
        705 : out = 27188;
        706 : out = 27132;
        707 : out = 27076;
        708 : out = 27019;
        709 : out = 26962;
        710 : out = 26905;
        711 : out = 26847;
        712 : out = 26789;
        713 : out = 26731;
        714 : out = 26673;
        715 : out = 26615;
        716 : out = 26556;
        717 : out = 26497;
        718 : out = 26437;
        719 : out = 26378;
        720 : out = 26318;
        721 : out = 26258;
        722 : out = 26198;
        723 : out = 26137;
        724 : out = 26077;
        725 : out = 26016;
        726 : out = 25954;
        727 : out = 25893;
        728 : out = 25831;
        729 : out = 25769;
        730 : out = 25707;
        731 : out = 25645;
        732 : out = 25582;
        733 : out = 25519;
        734 : out = 25456;
        735 : out = 25392;
        736 : out = 25329;
        737 : out = 25265;
        738 : out = 25201;
        739 : out = 25136;
        740 : out = 25072;
        741 : out = 25007;
        742 : out = 24942;
        743 : out = 24877;
        744 : out = 24811;
        745 : out = 24745;
        746 : out = 24679;
        747 : out = 24613;
        748 : out = 24546;
        749 : out = 24480;
        750 : out = 24413;
        751 : out = 24346;
        752 : out = 24278;
        753 : out = 24211;
        754 : out = 24143;
        755 : out = 24075;
        756 : out = 24006;
        757 : out = 23938;
        758 : out = 23869;
        759 : out = 23800;
        760 : out = 23731;
        761 : out = 23661;
        762 : out = 23592;
        763 : out = 23522;
        764 : out = 23452;
        765 : out = 23382;
        766 : out = 23311;
        767 : out = 23240;
        768 : out = 23169;
        769 : out = 23098;
        770 : out = 23027;
        771 : out = 22955;
        772 : out = 22883;
        773 : out = 22811;
        774 : out = 22739;
        775 : out = 22666;
        776 : out = 22594;
        777 : out = 22521;
        778 : out = 22448;
        779 : out = 22374;
        780 : out = 22301;
        781 : out = 22227;
        782 : out = 22153;
        783 : out = 22079;
        784 : out = 22004;
        785 : out = 21930;
        786 : out = 21855;
        787 : out = 21780;
        788 : out = 21705;
        789 : out = 21629;
        790 : out = 21554;
        791 : out = 21478;
        792 : out = 21402;
        793 : out = 21326;
        794 : out = 21249;
        795 : out = 21173;
        796 : out = 21096;
        797 : out = 21019;
        798 : out = 20942;
        799 : out = 20864;
        800 : out = 20787;
        801 : out = 20709;
        802 : out = 20631;
        803 : out = 20553;
        804 : out = 20474;
        805 : out = 20396;
        806 : out = 20317;
        807 : out = 20238;
        808 : out = 20159;
        809 : out = 20079;
        810 : out = 20000;
        811 : out = 19920;
        812 : out = 19840;
        813 : out = 19760;
        814 : out = 19680;
        815 : out = 19599;
        816 : out = 19519;
        817 : out = 19438;
        818 : out = 19357;
        819 : out = 19276;
        820 : out = 19194;
        821 : out = 19113;
        822 : out = 19031;
        823 : out = 18949;
        824 : out = 18867;
        825 : out = 18785;
        826 : out = 18702;
        827 : out = 18620;
        828 : out = 18537;
        829 : out = 18454;
        830 : out = 18371;
        831 : out = 18287;
        832 : out = 18204;
        833 : out = 18120;
        834 : out = 18036;
        835 : out = 17952;
        836 : out = 17868;
        837 : out = 17784;
        838 : out = 17699;
        839 : out = 17615;
        840 : out = 17530;
        841 : out = 17445;
        842 : out = 17360;
        843 : out = 17274;
        844 : out = 17189;
        845 : out = 17103;
        846 : out = 17017;
        847 : out = 16931;
        848 : out = 16845;
        849 : out = 16759;
        850 : out = 16672;
        851 : out = 16586;
        852 : out = 16499;
        853 : out = 16412;
        854 : out = 16325;
        855 : out = 16238;
        856 : out = 16150;
        857 : out = 16063;
        858 : out = 15975;
        859 : out = 15887;
        860 : out = 15799;
        861 : out = 15711;
        862 : out = 15623;
        863 : out = 15534;
        864 : out = 15446;
        865 : out = 15357;
        866 : out = 15268;
        867 : out = 15179;
        868 : out = 15090;
        869 : out = 15001;
        870 : out = 14911;
        871 : out = 14822;
        872 : out = 14732;
        873 : out = 14642;
        874 : out = 14552;
        875 : out = 14462;
        876 : out = 14372;
        877 : out = 14281;
        878 : out = 14191;
        879 : out = 14100;
        880 : out = 14009;
        881 : out = 13918;
        882 : out = 13827;
        883 : out = 13736;
        884 : out = 13645;
        885 : out = 13553;
        886 : out = 13462;
        887 : out = 13370;
        888 : out = 13278;
        889 : out = 13186;
        890 : out = 13094;
        891 : out = 13002;
        892 : out = 12909;
        893 : out = 12817;
        894 : out = 12724;
        895 : out = 12632;
        896 : out = 12539;
        897 : out = 12446;
        898 : out = 12353;
        899 : out = 12260;
        900 : out = 12166;
        901 : out = 12073;
        902 : out = 11980;
        903 : out = 11886;
        904 : out = 11792;
        905 : out = 11698;
        906 : out = 11604;
        907 : out = 11510;
        908 : out = 11416;
        909 : out = 11322;
        910 : out = 11227;
        911 : out = 11133;
        912 : out = 11038;
        913 : out = 10944;
        914 : out = 10849;
        915 : out = 10754;
        916 : out = 10659;
        917 : out = 10564;
        918 : out = 10469;
        919 : out = 10373;
        920 : out = 10278;
        921 : out = 10182;
        922 : out = 10087;
        923 : out = 9991;
        924 : out = 9895;
        925 : out = 9799;
        926 : out = 9703;
        927 : out = 9607;
        928 : out = 9511;
        929 : out = 9415;
        930 : out = 9319;
        931 : out = 9222;
        932 : out = 9126;
        933 : out = 9029;
        934 : out = 8932;
        935 : out = 8836;
        936 : out = 8739;
        937 : out = 8642;
        938 : out = 8545;
        939 : out = 8448;
        940 : out = 8351;
        941 : out = 8253;
        942 : out = 8156;
        943 : out = 8059;
        944 : out = 7961;
        945 : out = 7864;
        946 : out = 7766;
        947 : out = 7668;
        948 : out = 7571;
        949 : out = 7473;
        950 : out = 7375;
        951 : out = 7277;
        952 : out = 7179;
        953 : out = 7081;
        954 : out = 6982;
        955 : out = 6884;
        956 : out = 6786;
        957 : out = 6688;
        958 : out = 6589;
        959 : out = 6491;
        960 : out = 6392;
        961 : out = 6293;
        962 : out = 6195;
        963 : out = 6096;
        964 : out = 5997;
        965 : out = 5898;
        966 : out = 5799;
        967 : out = 5700;
        968 : out = 5601;
        969 : out = 5502;
        970 : out = 5403;
        971 : out = 5304;
        972 : out = 5205;
        973 : out = 5106;
        974 : out = 5006;
        975 : out = 4907;
        976 : out = 4807;
        977 : out = 4708;
        978 : out = 4608;
        979 : out = 4509;
        980 : out = 4409;
        981 : out = 4310;
        982 : out = 4210;
        983 : out = 4110;
        984 : out = 4011;
        985 : out = 3911;
        986 : out = 3811;
        987 : out = 3711;
        988 : out = 3611;
        989 : out = 3511;
        990 : out = 3411;
        991 : out = 3311;
        992 : out = 3211;
        993 : out = 3111;
        994 : out = 3011;
        995 : out = 2911;
        996 : out = 2811;
        997 : out = 2711;
        998 : out = 2610;
        999 : out = 2510;
        1000 : out = 2410;
        1001 : out = 2310;
        1002 : out = 2209;
        1003 : out = 2109;
        1004 : out = 2009;
        1005 : out = 1908;
        1006 : out = 1808;
        1007 : out = 1708;
        1008 : out = 1607;
        1009 : out = 1507;
        1010 : out = 1406;
        1011 : out = 1306;
        1012 : out = 1206;
        1013 : out = 1105;
        1014 : out = 1005;
        1015 : out = 904;
        1016 : out = 804;
        1017 : out = 703;
        1018 : out = 603;
        1019 : out = 502;
        1020 : out = 402;
        1021 : out = 301;
        1022 : out = 201;
        1023 : out = 100;
        1024 : out = 0;
        1025 : out = -100;
        1026 : out = -201;
        1027 : out = -301;
        1028 : out = -402;
        1029 : out = -502;
        1030 : out = -603;
        1031 : out = -703;
        1032 : out = -804;
        1033 : out = -904;
        1034 : out = -1005;
        1035 : out = -1105;
        1036 : out = -1206;
        1037 : out = -1306;
        1038 : out = -1406;
        1039 : out = -1507;
        1040 : out = -1607;
        1041 : out = -1708;
        1042 : out = -1808;
        1043 : out = -1908;
        1044 : out = -2009;
        1045 : out = -2109;
        1046 : out = -2209;
        1047 : out = -2310;
        1048 : out = -2410;
        1049 : out = -2510;
        1050 : out = -2610;
        1051 : out = -2711;
        1052 : out = -2811;
        1053 : out = -2911;
        1054 : out = -3011;
        1055 : out = -3111;
        1056 : out = -3211;
        1057 : out = -3311;
        1058 : out = -3411;
        1059 : out = -3511;
        1060 : out = -3611;
        1061 : out = -3711;
        1062 : out = -3811;
        1063 : out = -3911;
        1064 : out = -4011;
        1065 : out = -4110;
        1066 : out = -4210;
        1067 : out = -4310;
        1068 : out = -4409;
        1069 : out = -4509;
        1070 : out = -4608;
        1071 : out = -4708;
        1072 : out = -4807;
        1073 : out = -4907;
        1074 : out = -5006;
        1075 : out = -5106;
        1076 : out = -5205;
        1077 : out = -5304;
        1078 : out = -5403;
        1079 : out = -5502;
        1080 : out = -5601;
        1081 : out = -5700;
        1082 : out = -5799;
        1083 : out = -5898;
        1084 : out = -5997;
        1085 : out = -6096;
        1086 : out = -6195;
        1087 : out = -6293;
        1088 : out = -6392;
        1089 : out = -6491;
        1090 : out = -6589;
        1091 : out = -6688;
        1092 : out = -6786;
        1093 : out = -6884;
        1094 : out = -6982;
        1095 : out = -7081;
        1096 : out = -7179;
        1097 : out = -7277;
        1098 : out = -7375;
        1099 : out = -7473;
        1100 : out = -7571;
        1101 : out = -7668;
        1102 : out = -7766;
        1103 : out = -7864;
        1104 : out = -7961;
        1105 : out = -8059;
        1106 : out = -8156;
        1107 : out = -8253;
        1108 : out = -8351;
        1109 : out = -8448;
        1110 : out = -8545;
        1111 : out = -8642;
        1112 : out = -8739;
        1113 : out = -8836;
        1114 : out = -8932;
        1115 : out = -9029;
        1116 : out = -9126;
        1117 : out = -9222;
        1118 : out = -9319;
        1119 : out = -9415;
        1120 : out = -9511;
        1121 : out = -9607;
        1122 : out = -9703;
        1123 : out = -9799;
        1124 : out = -9895;
        1125 : out = -9991;
        1126 : out = -10087;
        1127 : out = -10182;
        1128 : out = -10278;
        1129 : out = -10373;
        1130 : out = -10469;
        1131 : out = -10564;
        1132 : out = -10659;
        1133 : out = -10754;
        1134 : out = -10849;
        1135 : out = -10944;
        1136 : out = -11038;
        1137 : out = -11133;
        1138 : out = -11227;
        1139 : out = -11322;
        1140 : out = -11416;
        1141 : out = -11510;
        1142 : out = -11604;
        1143 : out = -11698;
        1144 : out = -11792;
        1145 : out = -11886;
        1146 : out = -11980;
        1147 : out = -12073;
        1148 : out = -12166;
        1149 : out = -12260;
        1150 : out = -12353;
        1151 : out = -12446;
        1152 : out = -12539;
        1153 : out = -12632;
        1154 : out = -12724;
        1155 : out = -12817;
        1156 : out = -12909;
        1157 : out = -13002;
        1158 : out = -13094;
        1159 : out = -13186;
        1160 : out = -13278;
        1161 : out = -13370;
        1162 : out = -13462;
        1163 : out = -13553;
        1164 : out = -13645;
        1165 : out = -13736;
        1166 : out = -13827;
        1167 : out = -13918;
        1168 : out = -14009;
        1169 : out = -14100;
        1170 : out = -14191;
        1171 : out = -14281;
        1172 : out = -14372;
        1173 : out = -14462;
        1174 : out = -14552;
        1175 : out = -14642;
        1176 : out = -14732;
        1177 : out = -14822;
        1178 : out = -14911;
        1179 : out = -15001;
        1180 : out = -15090;
        1181 : out = -15179;
        1182 : out = -15268;
        1183 : out = -15357;
        1184 : out = -15446;
        1185 : out = -15534;
        1186 : out = -15623;
        1187 : out = -15711;
        1188 : out = -15799;
        1189 : out = -15887;
        1190 : out = -15975;
        1191 : out = -16063;
        1192 : out = -16150;
        1193 : out = -16238;
        1194 : out = -16325;
        1195 : out = -16412;
        1196 : out = -16499;
        1197 : out = -16586;
        1198 : out = -16672;
        1199 : out = -16759;
        1200 : out = -16845;
        1201 : out = -16931;
        1202 : out = -17017;
        1203 : out = -17103;
        1204 : out = -17189;
        1205 : out = -17274;
        1206 : out = -17360;
        1207 : out = -17445;
        1208 : out = -17530;
        1209 : out = -17615;
        1210 : out = -17699;
        1211 : out = -17784;
        1212 : out = -17868;
        1213 : out = -17952;
        1214 : out = -18036;
        1215 : out = -18120;
        1216 : out = -18204;
        1217 : out = -18287;
        1218 : out = -18371;
        1219 : out = -18454;
        1220 : out = -18537;
        1221 : out = -18620;
        1222 : out = -18702;
        1223 : out = -18785;
        1224 : out = -18867;
        1225 : out = -18949;
        1226 : out = -19031;
        1227 : out = -19113;
        1228 : out = -19194;
        1229 : out = -19276;
        1230 : out = -19357;
        1231 : out = -19438;
        1232 : out = -19519;
        1233 : out = -19599;
        1234 : out = -19680;
        1235 : out = -19760;
        1236 : out = -19840;
        1237 : out = -19920;
        1238 : out = -20000;
        1239 : out = -20079;
        1240 : out = -20159;
        1241 : out = -20238;
        1242 : out = -20317;
        1243 : out = -20396;
        1244 : out = -20474;
        1245 : out = -20553;
        1246 : out = -20631;
        1247 : out = -20709;
        1248 : out = -20787;
        1249 : out = -20864;
        1250 : out = -20942;
        1251 : out = -21019;
        1252 : out = -21096;
        1253 : out = -21173;
        1254 : out = -21249;
        1255 : out = -21326;
        1256 : out = -21402;
        1257 : out = -21478;
        1258 : out = -21554;
        1259 : out = -21629;
        1260 : out = -21705;
        1261 : out = -21780;
        1262 : out = -21855;
        1263 : out = -21930;
        1264 : out = -22004;
        1265 : out = -22079;
        1266 : out = -22153;
        1267 : out = -22227;
        1268 : out = -22301;
        1269 : out = -22374;
        1270 : out = -22448;
        1271 : out = -22521;
        1272 : out = -22594;
        1273 : out = -22666;
        1274 : out = -22739;
        1275 : out = -22811;
        1276 : out = -22883;
        1277 : out = -22955;
        1278 : out = -23027;
        1279 : out = -23098;
        1280 : out = -23169;
        1281 : out = -23240;
        1282 : out = -23311;
        1283 : out = -23382;
        1284 : out = -23452;
        1285 : out = -23522;
        1286 : out = -23592;
        1287 : out = -23661;
        1288 : out = -23731;
        1289 : out = -23800;
        1290 : out = -23869;
        1291 : out = -23938;
        1292 : out = -24006;
        1293 : out = -24075;
        1294 : out = -24143;
        1295 : out = -24211;
        1296 : out = -24278;
        1297 : out = -24346;
        1298 : out = -24413;
        1299 : out = -24480;
        1300 : out = -24546;
        1301 : out = -24613;
        1302 : out = -24679;
        1303 : out = -24745;
        1304 : out = -24811;
        1305 : out = -24877;
        1306 : out = -24942;
        1307 : out = -25007;
        1308 : out = -25072;
        1309 : out = -25136;
        1310 : out = -25201;
        1311 : out = -25265;
        1312 : out = -25329;
        1313 : out = -25392;
        1314 : out = -25456;
        1315 : out = -25519;
        1316 : out = -25582;
        1317 : out = -25645;
        1318 : out = -25707;
        1319 : out = -25769;
        1320 : out = -25831;
        1321 : out = -25893;
        1322 : out = -25954;
        1323 : out = -26016;
        1324 : out = -26077;
        1325 : out = -26137;
        1326 : out = -26198;
        1327 : out = -26258;
        1328 : out = -26318;
        1329 : out = -26378;
        1330 : out = -26437;
        1331 : out = -26497;
        1332 : out = -26556;
        1333 : out = -26615;
        1334 : out = -26673;
        1335 : out = -26731;
        1336 : out = -26789;
        1337 : out = -26847;
        1338 : out = -26905;
        1339 : out = -26962;
        1340 : out = -27019;
        1341 : out = -27076;
        1342 : out = -27132;
        1343 : out = -27188;
        1344 : out = -27244;
        1345 : out = -27300;
        1346 : out = -27355;
        1347 : out = -27411;
        1348 : out = -27466;
        1349 : out = -27520;
        1350 : out = -27575;
        1351 : out = -27629;
        1352 : out = -27683;
        1353 : out = -27736;
        1354 : out = -27790;
        1355 : out = -27843;
        1356 : out = -27896;
        1357 : out = -27948;
        1358 : out = -28001;
        1359 : out = -28053;
        1360 : out = -28105;
        1361 : out = -28156;
        1362 : out = -28208;
        1363 : out = -28259;
        1364 : out = -28309;
        1365 : out = -28360;
        1366 : out = -28410;
        1367 : out = -28460;
        1368 : out = -28510;
        1369 : out = -28559;
        1370 : out = -28608;
        1371 : out = -28657;
        1372 : out = -28706;
        1373 : out = -28754;
        1374 : out = -28802;
        1375 : out = -28850;
        1376 : out = -28897;
        1377 : out = -28945;
        1378 : out = -28992;
        1379 : out = -29038;
        1380 : out = -29085;
        1381 : out = -29131;
        1382 : out = -29177;
        1383 : out = -29222;
        1384 : out = -29268;
        1385 : out = -29313;
        1386 : out = -29358;
        1387 : out = -29402;
        1388 : out = -29446;
        1389 : out = -29490;
        1390 : out = -29534;
        1391 : out = -29577;
        1392 : out = -29621;
        1393 : out = -29663;
        1394 : out = -29706;
        1395 : out = -29748;
        1396 : out = -29790;
        1397 : out = -29832;
        1398 : out = -29873;
        1399 : out = -29915;
        1400 : out = -29955;
        1401 : out = -29996;
        1402 : out = -30036;
        1403 : out = -30076;
        1404 : out = -30116;
        1405 : out = -30156;
        1406 : out = -30195;
        1407 : out = -30234;
        1408 : out = -30272;
        1409 : out = -30311;
        1410 : out = -30349;
        1411 : out = -30386;
        1412 : out = -30424;
        1413 : out = -30461;
        1414 : out = -30498;
        1415 : out = -30535;
        1416 : out = -30571;
        1417 : out = -30607;
        1418 : out = -30643;
        1419 : out = -30678;
        1420 : out = -30713;
        1421 : out = -30748;
        1422 : out = -30783;
        1423 : out = -30817;
        1424 : out = -30851;
        1425 : out = -30885;
        1426 : out = -30918;
        1427 : out = -30951;
        1428 : out = -30984;
        1429 : out = -31017;
        1430 : out = -31049;
        1431 : out = -31081;
        1432 : out = -31113;
        1433 : out = -31144;
        1434 : out = -31175;
        1435 : out = -31206;
        1436 : out = -31236;
        1437 : out = -31267;
        1438 : out = -31297;
        1439 : out = -31326;
        1440 : out = -31356;
        1441 : out = -31385;
        1442 : out = -31413;
        1443 : out = -31442;
        1444 : out = -31470;
        1445 : out = -31498;
        1446 : out = -31525;
        1447 : out = -31553;
        1448 : out = -31580;
        1449 : out = -31606;
        1450 : out = -31633;
        1451 : out = -31659;
        1452 : out = -31684;
        1453 : out = -31710;
        1454 : out = -31735;
        1455 : out = -31760;
        1456 : out = -31785;
        1457 : out = -31809;
        1458 : out = -31833;
        1459 : out = -31856;
        1460 : out = -31880;
        1461 : out = -31903;
        1462 : out = -31926;
        1463 : out = -31948;
        1464 : out = -31970;
        1465 : out = -31992;
        1466 : out = -32014;
        1467 : out = -32035;
        1468 : out = -32056;
        1469 : out = -32077;
        1470 : out = -32097;
        1471 : out = -32117;
        1472 : out = -32137;
        1473 : out = -32156;
        1474 : out = -32176;
        1475 : out = -32194;
        1476 : out = -32213;
        1477 : out = -32231;
        1478 : out = -32249;
        1479 : out = -32267;
        1480 : out = -32284;
        1481 : out = -32301;
        1482 : out = -32318;
        1483 : out = -32334;
        1484 : out = -32350;
        1485 : out = -32366;
        1486 : out = -32382;
        1487 : out = -32397;
        1488 : out = -32412;
        1489 : out = -32426;
        1490 : out = -32441;
        1491 : out = -32455;
        1492 : out = -32468;
        1493 : out = -32482;
        1494 : out = -32495;
        1495 : out = -32508;
        1496 : out = -32520;
        1497 : out = -32532;
        1498 : out = -32544;
        1499 : out = -32556;
        1500 : out = -32567;
        1501 : out = -32578;
        1502 : out = -32588;
        1503 : out = -32599;
        1504 : out = -32609;
        1505 : out = -32618;
        1506 : out = -32628;
        1507 : out = -32637;
        1508 : out = -32646;
        1509 : out = -32654;
        1510 : out = -32662;
        1511 : out = -32670;
        1512 : out = -32678;
        1513 : out = -32685;
        1514 : out = -32692;
        1515 : out = -32699;
        1516 : out = -32705;
        1517 : out = -32711;
        1518 : out = -32717;
        1519 : out = -32722;
        1520 : out = -32727;
        1521 : out = -32732;
        1522 : out = -32736;
        1523 : out = -32740;
        1524 : out = -32744;
        1525 : out = -32748;
        1526 : out = -32751;
        1527 : out = -32754;
        1528 : out = -32757;
        1529 : out = -32759;
        1530 : out = -32761;
        1531 : out = -32763;
        1532 : out = -32764;
        1533 : out = -32765;
        1534 : out = -32766;
        1535 : out = -32766;
        1536 : out = -32767;
        1537 : out = -32766;
        1538 : out = -32766;
        1539 : out = -32765;
        1540 : out = -32764;
        1541 : out = -32763;
        1542 : out = -32761;
        1543 : out = -32759;
        1544 : out = -32757;
        1545 : out = -32754;
        1546 : out = -32751;
        1547 : out = -32748;
        1548 : out = -32744;
        1549 : out = -32740;
        1550 : out = -32736;
        1551 : out = -32732;
        1552 : out = -32727;
        1553 : out = -32722;
        1554 : out = -32717;
        1555 : out = -32711;
        1556 : out = -32705;
        1557 : out = -32699;
        1558 : out = -32692;
        1559 : out = -32685;
        1560 : out = -32678;
        1561 : out = -32670;
        1562 : out = -32662;
        1563 : out = -32654;
        1564 : out = -32646;
        1565 : out = -32637;
        1566 : out = -32628;
        1567 : out = -32618;
        1568 : out = -32609;
        1569 : out = -32599;
        1570 : out = -32588;
        1571 : out = -32578;
        1572 : out = -32567;
        1573 : out = -32556;
        1574 : out = -32544;
        1575 : out = -32532;
        1576 : out = -32520;
        1577 : out = -32508;
        1578 : out = -32495;
        1579 : out = -32482;
        1580 : out = -32468;
        1581 : out = -32455;
        1582 : out = -32441;
        1583 : out = -32426;
        1584 : out = -32412;
        1585 : out = -32397;
        1586 : out = -32382;
        1587 : out = -32366;
        1588 : out = -32350;
        1589 : out = -32334;
        1590 : out = -32318;
        1591 : out = -32301;
        1592 : out = -32284;
        1593 : out = -32267;
        1594 : out = -32249;
        1595 : out = -32231;
        1596 : out = -32213;
        1597 : out = -32194;
        1598 : out = -32176;
        1599 : out = -32156;
        1600 : out = -32137;
        1601 : out = -32117;
        1602 : out = -32097;
        1603 : out = -32077;
        1604 : out = -32056;
        1605 : out = -32035;
        1606 : out = -32014;
        1607 : out = -31992;
        1608 : out = -31970;
        1609 : out = -31948;
        1610 : out = -31926;
        1611 : out = -31903;
        1612 : out = -31880;
        1613 : out = -31856;
        1614 : out = -31833;
        1615 : out = -31809;
        1616 : out = -31785;
        1617 : out = -31760;
        1618 : out = -31735;
        1619 : out = -31710;
        1620 : out = -31684;
        1621 : out = -31659;
        1622 : out = -31633;
        1623 : out = -31606;
        1624 : out = -31580;
        1625 : out = -31553;
        1626 : out = -31525;
        1627 : out = -31498;
        1628 : out = -31470;
        1629 : out = -31442;
        1630 : out = -31413;
        1631 : out = -31385;
        1632 : out = -31356;
        1633 : out = -31326;
        1634 : out = -31297;
        1635 : out = -31267;
        1636 : out = -31236;
        1637 : out = -31206;
        1638 : out = -31175;
        1639 : out = -31144;
        1640 : out = -31113;
        1641 : out = -31081;
        1642 : out = -31049;
        1643 : out = -31017;
        1644 : out = -30984;
        1645 : out = -30951;
        1646 : out = -30918;
        1647 : out = -30885;
        1648 : out = -30851;
        1649 : out = -30817;
        1650 : out = -30783;
        1651 : out = -30748;
        1652 : out = -30713;
        1653 : out = -30678;
        1654 : out = -30643;
        1655 : out = -30607;
        1656 : out = -30571;
        1657 : out = -30535;
        1658 : out = -30498;
        1659 : out = -30461;
        1660 : out = -30424;
        1661 : out = -30386;
        1662 : out = -30349;
        1663 : out = -30311;
        1664 : out = -30272;
        1665 : out = -30234;
        1666 : out = -30195;
        1667 : out = -30156;
        1668 : out = -30116;
        1669 : out = -30076;
        1670 : out = -30036;
        1671 : out = -29996;
        1672 : out = -29955;
        1673 : out = -29915;
        1674 : out = -29873;
        1675 : out = -29832;
        1676 : out = -29790;
        1677 : out = -29748;
        1678 : out = -29706;
        1679 : out = -29663;
        1680 : out = -29621;
        1681 : out = -29577;
        1682 : out = -29534;
        1683 : out = -29490;
        1684 : out = -29446;
        1685 : out = -29402;
        1686 : out = -29358;
        1687 : out = -29313;
        1688 : out = -29268;
        1689 : out = -29222;
        1690 : out = -29177;
        1691 : out = -29131;
        1692 : out = -29085;
        1693 : out = -29038;
        1694 : out = -28992;
        1695 : out = -28945;
        1696 : out = -28897;
        1697 : out = -28850;
        1698 : out = -28802;
        1699 : out = -28754;
        1700 : out = -28706;
        1701 : out = -28657;
        1702 : out = -28608;
        1703 : out = -28559;
        1704 : out = -28510;
        1705 : out = -28460;
        1706 : out = -28410;
        1707 : out = -28360;
        1708 : out = -28309;
        1709 : out = -28259;
        1710 : out = -28208;
        1711 : out = -28156;
        1712 : out = -28105;
        1713 : out = -28053;
        1714 : out = -28001;
        1715 : out = -27948;
        1716 : out = -27896;
        1717 : out = -27843;
        1718 : out = -27790;
        1719 : out = -27736;
        1720 : out = -27683;
        1721 : out = -27629;
        1722 : out = -27575;
        1723 : out = -27520;
        1724 : out = -27466;
        1725 : out = -27411;
        1726 : out = -27355;
        1727 : out = -27300;
        1728 : out = -27244;
        1729 : out = -27188;
        1730 : out = -27132;
        1731 : out = -27076;
        1732 : out = -27019;
        1733 : out = -26962;
        1734 : out = -26905;
        1735 : out = -26847;
        1736 : out = -26789;
        1737 : out = -26731;
        1738 : out = -26673;
        1739 : out = -26615;
        1740 : out = -26556;
        1741 : out = -26497;
        1742 : out = -26437;
        1743 : out = -26378;
        1744 : out = -26318;
        1745 : out = -26258;
        1746 : out = -26198;
        1747 : out = -26137;
        1748 : out = -26077;
        1749 : out = -26016;
        1750 : out = -25954;
        1751 : out = -25893;
        1752 : out = -25831;
        1753 : out = -25769;
        1754 : out = -25707;
        1755 : out = -25645;
        1756 : out = -25582;
        1757 : out = -25519;
        1758 : out = -25456;
        1759 : out = -25392;
        1760 : out = -25329;
        1761 : out = -25265;
        1762 : out = -25201;
        1763 : out = -25136;
        1764 : out = -25072;
        1765 : out = -25007;
        1766 : out = -24942;
        1767 : out = -24877;
        1768 : out = -24811;
        1769 : out = -24745;
        1770 : out = -24679;
        1771 : out = -24613;
        1772 : out = -24546;
        1773 : out = -24480;
        1774 : out = -24413;
        1775 : out = -24346;
        1776 : out = -24278;
        1777 : out = -24211;
        1778 : out = -24143;
        1779 : out = -24075;
        1780 : out = -24006;
        1781 : out = -23938;
        1782 : out = -23869;
        1783 : out = -23800;
        1784 : out = -23731;
        1785 : out = -23661;
        1786 : out = -23592;
        1787 : out = -23522;
        1788 : out = -23452;
        1789 : out = -23382;
        1790 : out = -23311;
        1791 : out = -23240;
        1792 : out = -23169;
        1793 : out = -23098;
        1794 : out = -23027;
        1795 : out = -22955;
        1796 : out = -22883;
        1797 : out = -22811;
        1798 : out = -22739;
        1799 : out = -22666;
        1800 : out = -22594;
        1801 : out = -22521;
        1802 : out = -22448;
        1803 : out = -22374;
        1804 : out = -22301;
        1805 : out = -22227;
        1806 : out = -22153;
        1807 : out = -22079;
        1808 : out = -22004;
        1809 : out = -21930;
        1810 : out = -21855;
        1811 : out = -21780;
        1812 : out = -21705;
        1813 : out = -21629;
        1814 : out = -21554;
        1815 : out = -21478;
        1816 : out = -21402;
        1817 : out = -21326;
        1818 : out = -21249;
        1819 : out = -21173;
        1820 : out = -21096;
        1821 : out = -21019;
        1822 : out = -20942;
        1823 : out = -20864;
        1824 : out = -20787;
        1825 : out = -20709;
        1826 : out = -20631;
        1827 : out = -20553;
        1828 : out = -20474;
        1829 : out = -20396;
        1830 : out = -20317;
        1831 : out = -20238;
        1832 : out = -20159;
        1833 : out = -20079;
        1834 : out = -20000;
        1835 : out = -19920;
        1836 : out = -19840;
        1837 : out = -19760;
        1838 : out = -19680;
        1839 : out = -19599;
        1840 : out = -19519;
        1841 : out = -19438;
        1842 : out = -19357;
        1843 : out = -19276;
        1844 : out = -19194;
        1845 : out = -19113;
        1846 : out = -19031;
        1847 : out = -18949;
        1848 : out = -18867;
        1849 : out = -18785;
        1850 : out = -18702;
        1851 : out = -18620;
        1852 : out = -18537;
        1853 : out = -18454;
        1854 : out = -18371;
        1855 : out = -18287;
        1856 : out = -18204;
        1857 : out = -18120;
        1858 : out = -18036;
        1859 : out = -17952;
        1860 : out = -17868;
        1861 : out = -17784;
        1862 : out = -17699;
        1863 : out = -17615;
        1864 : out = -17530;
        1865 : out = -17445;
        1866 : out = -17360;
        1867 : out = -17274;
        1868 : out = -17189;
        1869 : out = -17103;
        1870 : out = -17017;
        1871 : out = -16931;
        1872 : out = -16845;
        1873 : out = -16759;
        1874 : out = -16672;
        1875 : out = -16586;
        1876 : out = -16499;
        1877 : out = -16412;
        1878 : out = -16325;
        1879 : out = -16238;
        1880 : out = -16150;
        1881 : out = -16063;
        1882 : out = -15975;
        1883 : out = -15887;
        1884 : out = -15799;
        1885 : out = -15711;
        1886 : out = -15623;
        1887 : out = -15534;
        1888 : out = -15446;
        1889 : out = -15357;
        1890 : out = -15268;
        1891 : out = -15179;
        1892 : out = -15090;
        1893 : out = -15001;
        1894 : out = -14911;
        1895 : out = -14822;
        1896 : out = -14732;
        1897 : out = -14642;
        1898 : out = -14552;
        1899 : out = -14462;
        1900 : out = -14372;
        1901 : out = -14281;
        1902 : out = -14191;
        1903 : out = -14100;
        1904 : out = -14009;
        1905 : out = -13918;
        1906 : out = -13827;
        1907 : out = -13736;
        1908 : out = -13645;
        1909 : out = -13553;
        1910 : out = -13462;
        1911 : out = -13370;
        1912 : out = -13278;
        1913 : out = -13186;
        1914 : out = -13094;
        1915 : out = -13002;
        1916 : out = -12909;
        1917 : out = -12817;
        1918 : out = -12724;
        1919 : out = -12632;
        1920 : out = -12539;
        1921 : out = -12446;
        1922 : out = -12353;
        1923 : out = -12260;
        1924 : out = -12166;
        1925 : out = -12073;
        1926 : out = -11980;
        1927 : out = -11886;
        1928 : out = -11792;
        1929 : out = -11698;
        1930 : out = -11604;
        1931 : out = -11510;
        1932 : out = -11416;
        1933 : out = -11322;
        1934 : out = -11227;
        1935 : out = -11133;
        1936 : out = -11038;
        1937 : out = -10944;
        1938 : out = -10849;
        1939 : out = -10754;
        1940 : out = -10659;
        1941 : out = -10564;
        1942 : out = -10469;
        1943 : out = -10373;
        1944 : out = -10278;
        1945 : out = -10182;
        1946 : out = -10087;
        1947 : out = -9991;
        1948 : out = -9895;
        1949 : out = -9799;
        1950 : out = -9703;
        1951 : out = -9607;
        1952 : out = -9511;
        1953 : out = -9415;
        1954 : out = -9319;
        1955 : out = -9222;
        1956 : out = -9126;
        1957 : out = -9029;
        1958 : out = -8932;
        1959 : out = -8836;
        1960 : out = -8739;
        1961 : out = -8642;
        1962 : out = -8545;
        1963 : out = -8448;
        1964 : out = -8351;
        1965 : out = -8253;
        1966 : out = -8156;
        1967 : out = -8059;
        1968 : out = -7961;
        1969 : out = -7864;
        1970 : out = -7766;
        1971 : out = -7668;
        1972 : out = -7571;
        1973 : out = -7473;
        1974 : out = -7375;
        1975 : out = -7277;
        1976 : out = -7179;
        1977 : out = -7081;
        1978 : out = -6982;
        1979 : out = -6884;
        1980 : out = -6786;
        1981 : out = -6688;
        1982 : out = -6589;
        1983 : out = -6491;
        1984 : out = -6392;
        1985 : out = -6293;
        1986 : out = -6195;
        1987 : out = -6096;
        1988 : out = -5997;
        1989 : out = -5898;
        1990 : out = -5799;
        1991 : out = -5700;
        1992 : out = -5601;
        1993 : out = -5502;
        1994 : out = -5403;
        1995 : out = -5304;
        1996 : out = -5205;
        1997 : out = -5106;
        1998 : out = -5006;
        1999 : out = -4907;
        2000 : out = -4807;
        2001 : out = -4708;
        2002 : out = -4608;
        2003 : out = -4509;
        2004 : out = -4409;
        2005 : out = -4310;
        2006 : out = -4210;
        2007 : out = -4110;
        2008 : out = -4011;
        2009 : out = -3911;
        2010 : out = -3811;
        2011 : out = -3711;
        2012 : out = -3611;
        2013 : out = -3511;
        2014 : out = -3411;
        2015 : out = -3311;
        2016 : out = -3211;
        2017 : out = -3111;
        2018 : out = -3011;
        2019 : out = -2911;
        2020 : out = -2811;
        2021 : out = -2711;
        2022 : out = -2610;
        2023 : out = -2510;
        2024 : out = -2410;
        2025 : out = -2310;
        2026 : out = -2209;
        2027 : out = -2109;
        2028 : out = -2009;
        2029 : out = -1908;
        2030 : out = -1808;
        2031 : out = -1708;
        2032 : out = -1607;
        2033 : out = -1507;
        2034 : out = -1406;
        2035 : out = -1306;
        2036 : out = -1206;
        2037 : out = -1105;
        2038 : out = -1005;
        2039 : out = -904;
        2040 : out = -804;
        2041 : out = -703;
        2042 : out = -603;
        2043 : out = -502;
        2044 : out = -402;
        2045 : out = -301;
        2046 : out = -201;
        2047 : out = -100;
    endcase
end
endmodule
