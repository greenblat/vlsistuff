module exptab ( input [9:0] index,output [31:0] result);
assign result = 
    (index==0) ? 32'h40000000 : 
    (index==1) ? 32'h40001630 : 
    (index==2) ? 32'h40002c64 : 
    (index==3) ? 32'h4000429c : 
    (index==4) ? 32'h400058d7 : 
    (index==5) ? 32'h40006f17 : 
    (index==6) ? 32'h4000855a : 
    (index==7) ? 32'h40009ba2 : 
    (index==8) ? 32'h4000b1ed : 
    (index==9) ? 32'h4000c83c : 
    (index==10) ? 32'h4000de8f : 
    (index==11) ? 32'h4000f4e5 : 
    (index==12) ? 32'h40010b40 : 
    (index==13) ? 32'h4001219f : 
    (index==14) ? 32'h40013801 : 
    (index==15) ? 32'h40014e67 : 
    (index==16) ? 32'h400164d1 : 
    (index==17) ? 32'h40017b3f : 
    (index==18) ? 32'h400191b1 : 
    (index==19) ? 32'h4001a827 : 
    (index==20) ? 32'h4001bea1 : 
    (index==21) ? 32'h4001d51f : 
    (index==22) ? 32'h4001eba0 : 
    (index==23) ? 32'h40020225 : 
    (index==24) ? 32'h400218af : 
    (index==25) ? 32'h40022f3c : 
    (index==26) ? 32'h400245cd : 
    (index==27) ? 32'h40025c62 : 
    (index==28) ? 32'h400272fb : 
    (index==29) ? 32'h40028998 : 
    (index==30) ? 32'h4002a039 : 
    (index==31) ? 32'h4002b6dd : 
    (index==32) ? 32'h4002cd86 : 
    (index==33) ? 32'h4002e433 : 
    (index==34) ? 32'h4002fae3 : 
    (index==35) ? 32'h40031198 : 
    (index==36) ? 32'h40032850 : 
    (index==37) ? 32'h40033f0c : 
    (index==38) ? 32'h400355cc : 
    (index==39) ? 32'h40036c91 : 
    (index==40) ? 32'h40038359 : 
    (index==41) ? 32'h40039a25 : 
    (index==42) ? 32'h4003b0f5 : 
    (index==43) ? 32'h4003c7c9 : 
    (index==44) ? 32'h4003dea1 : 
    (index==45) ? 32'h4003f57d : 
    (index==46) ? 32'h40040c5d : 
    (index==47) ? 32'h40042340 : 
    (index==48) ? 32'h40043a28 : 
    (index==49) ? 32'h40045114 : 
    (index==50) ? 32'h40046804 : 
    (index==51) ? 32'h40047ef8 : 
    (index==52) ? 32'h400495ef : 
    (index==53) ? 32'h4004aceb : 
    (index==54) ? 32'h4004c3eb : 
    (index==55) ? 32'h4004daee : 
    (index==56) ? 32'h4004f1f6 : 
    (index==57) ? 32'h40050901 : 
    (index==58) ? 32'h40052011 : 
    (index==59) ? 32'h40053725 : 
    (index==60) ? 32'h40054e3c : 
    (index==61) ? 32'h40056558 : 
    (index==62) ? 32'h40057c78 : 
    (index==63) ? 32'h4005939b : 
    (index==64) ? 32'h4005aac3 : 
    (index==65) ? 32'h4005c1ef : 
    (index==66) ? 32'h4005d91e : 
    (index==67) ? 32'h4005f052 : 
    (index==68) ? 32'h4006078a : 
    (index==69) ? 32'h40061ec5 : 
    (index==70) ? 32'h40063605 : 
    (index==71) ? 32'h40064d49 : 
    (index==72) ? 32'h40066491 : 
    (index==73) ? 32'h40067bdd : 
    (index==74) ? 32'h4006932d : 
    (index==75) ? 32'h4006aa81 : 
    (index==76) ? 32'h4006c1d9 : 
    (index==77) ? 32'h4006d935 : 
    (index==78) ? 32'h4006f095 : 
    (index==79) ? 32'h400707f9 : 
    (index==80) ? 32'h40071f61 : 
    (index==81) ? 32'h400736cd : 
    (index==82) ? 32'h40074e3e : 
    (index==83) ? 32'h400765b2 : 
    (index==84) ? 32'h40077d2a : 
    (index==85) ? 32'h400794a7 : 
    (index==86) ? 32'h4007ac28 : 
    (index==87) ? 32'h4007c3ac : 
    (index==88) ? 32'h4007db35 : 
    (index==89) ? 32'h4007f2c2 : 
    (index==90) ? 32'h40080a53 : 
    (index==91) ? 32'h400821e8 : 
    (index==92) ? 32'h40083981 : 
    (index==93) ? 32'h4008511e : 
    (index==94) ? 32'h400868bf : 
    (index==95) ? 32'h40088065 : 
    (index==96) ? 32'h4008980e : 
    (index==97) ? 32'h4008afbc : 
    (index==98) ? 32'h4008c76d : 
    (index==99) ? 32'h4008df23 : 
    (index==100) ? 32'h4008f6dd : 
    (index==101) ? 32'h40090e9b : 
    (index==102) ? 32'h4009265d : 
    (index==103) ? 32'h40093e23 : 
    (index==104) ? 32'h400955ee : 
    (index==105) ? 32'h40096dbc : 
    (index==106) ? 32'h4009858f : 
    (index==107) ? 32'h40099d65 : 
    (index==108) ? 32'h4009b540 : 
    (index==109) ? 32'h4009cd1f : 
    (index==110) ? 32'h4009e502 : 
    (index==111) ? 32'h4009fcea : 
    (index==112) ? 32'h400a14d5 : 
    (index==113) ? 32'h400a2cc5 : 
    (index==114) ? 32'h400a44b8 : 
    (index==115) ? 32'h400a5cb0 : 
    (index==116) ? 32'h400a74ac : 
    (index==117) ? 32'h400a8cac : 
    (index==118) ? 32'h400aa4b1 : 
    (index==119) ? 32'h400abcb9 : 
    (index==120) ? 32'h400ad4c6 : 
    (index==121) ? 32'h400aecd7 : 
    (index==122) ? 32'h400b04ec : 
    (index==123) ? 32'h400b1d05 : 
    (index==124) ? 32'h400b3522 : 
    (index==125) ? 32'h400b4d44 : 
    (index==126) ? 32'h400b6569 : 
    (index==127) ? 32'h400b7d93 : 
    (index==128) ? 32'h400b95c1 : 
    (index==129) ? 32'h400badf4 : 
    (index==130) ? 32'h400bc62a : 
    (index==131) ? 32'h400bde65 : 
    (index==132) ? 32'h400bf6a4 : 
    (index==133) ? 32'h400c0ee7 : 
    (index==134) ? 32'h400c272e : 
    (index==135) ? 32'h400c3f7a : 
    (index==136) ? 32'h400c57c9 : 
    (index==137) ? 32'h400c701d : 
    (index==138) ? 32'h400c8875 : 
    (index==139) ? 32'h400ca0d2 : 
    (index==140) ? 32'h400cb932 : 
    (index==141) ? 32'h400cd197 : 
    (index==142) ? 32'h400cea00 : 
    (index==143) ? 32'h400d026d : 
    (index==144) ? 32'h400d1adf : 
    (index==145) ? 32'h400d3355 : 
    (index==146) ? 32'h400d4bcf : 
    (index==147) ? 32'h400d644d : 
    (index==148) ? 32'h400d7ccf : 
    (index==149) ? 32'h400d9556 : 
    (index==150) ? 32'h400dade1 : 
    (index==151) ? 32'h400dc670 : 
    (index==152) ? 32'h400ddf04 : 
    (index==153) ? 32'h400df79b : 
    (index==154) ? 32'h400e1037 : 
    (index==155) ? 32'h400e28d8 : 
    (index==156) ? 32'h400e417c : 
    (index==157) ? 32'h400e5a25 : 
    (index==158) ? 32'h400e72d2 : 
    (index==159) ? 32'h400e8b83 : 
    (index==160) ? 32'h400ea439 : 
    (index==161) ? 32'h400ebcf3 : 
    (index==162) ? 32'h400ed5b1 : 
    (index==163) ? 32'h400eee74 : 
    (index==164) ? 32'h400f073a : 
    (index==165) ? 32'h400f2006 : 
    (index==166) ? 32'h400f38d5 : 
    (index==167) ? 32'h400f51a9 : 
    (index==168) ? 32'h400f6a81 : 
    (index==169) ? 32'h400f835d : 
    (index==170) ? 32'h400f9c3d : 
    (index==171) ? 32'h400fb522 : 
    (index==172) ? 32'h400fce0c : 
    (index==173) ? 32'h400fe6f9 : 
    (index==174) ? 32'h400fffeb : 
    (index==175) ? 32'h401018e1 : 
    (index==176) ? 32'h401031dc : 
    (index==177) ? 32'h40104adb : 
    (index==178) ? 32'h401063de : 
    (index==179) ? 32'h40107ce5 : 
    (index==180) ? 32'h401095f1 : 
    (index==181) ? 32'h4010af01 : 
    (index==182) ? 32'h4010c816 : 
    (index==183) ? 32'h4010e12f : 
    (index==184) ? 32'h4010fa4c : 
    (index==185) ? 32'h4011136e : 
    (index==186) ? 32'h40112c94 : 
    (index==187) ? 32'h401145be : 
    (index==188) ? 32'h40115eed : 
    (index==189) ? 32'h40117820 : 
    (index==190) ? 32'h40119157 : 
    (index==191) ? 32'h4011aa93 : 
    (index==192) ? 32'h4011c3d3 : 
    (index==193) ? 32'h4011dd17 : 
    (index==194) ? 32'h4011f660 : 
    (index==195) ? 32'h40120fae : 
    (index==196) ? 32'h401228ff : 
    (index==197) ? 32'h40124255 : 
    (index==198) ? 32'h40125bb0 : 
    (index==199) ? 32'h4012750f : 
    (index==200) ? 32'h40128e72 : 
    (index==201) ? 32'h4012a7da : 
    (index==202) ? 32'h4012c146 : 
    (index==203) ? 32'h4012dab6 : 
    (index==204) ? 32'h4012f42b : 
    (index==205) ? 32'h40130da4 : 
    (index==206) ? 32'h40132722 : 
    (index==207) ? 32'h401340a4 : 
    (index==208) ? 32'h40135a2b : 
    (index==209) ? 32'h401373b6 : 
    (index==210) ? 32'h40138d45 : 
    (index==211) ? 32'h4013a6d9 : 
    (index==212) ? 32'h4013c071 : 
    (index==213) ? 32'h4013da0e : 
    (index==214) ? 32'h4013f3af : 
    (index==215) ? 32'h40140d55 : 
    (index==216) ? 32'h401426ff : 
    (index==217) ? 32'h401440ad : 
    (index==218) ? 32'h40145a60 : 
    (index==219) ? 32'h40147417 : 
    (index==220) ? 32'h40148dd3 : 
    (index==221) ? 32'h4014a793 : 
    (index==222) ? 32'h4014c158 : 
    (index==223) ? 32'h4014db21 : 
    (index==224) ? 32'h4014f4ef : 
    (index==225) ? 32'h40150ec1 : 
    (index==226) ? 32'h40152898 : 
    (index==227) ? 32'h40154273 : 
    (index==228) ? 32'h40155c53 : 
    (index==229) ? 32'h40157637 : 
    (index==230) ? 32'h4015901f : 
    (index==231) ? 32'h4015aa0c : 
    (index==232) ? 32'h4015c3fe : 
    (index==233) ? 32'h4015ddf4 : 
    (index==234) ? 32'h4015f7ef : 
    (index==235) ? 32'h401611ee : 
    (index==236) ? 32'h40162bf1 : 
    (index==237) ? 32'h401645f9 : 
    (index==238) ? 32'h40166006 : 
    (index==239) ? 32'h40167a17 : 
    (index==240) ? 32'h4016942d : 
    (index==241) ? 32'h4016ae47 : 
    (index==242) ? 32'h4016c866 : 
    (index==243) ? 32'h4016e289 : 
    (index==244) ? 32'h4016fcb0 : 
    (index==245) ? 32'h401716dd : 
    (index==246) ? 32'h4017310e : 
    (index==247) ? 32'h40174b43 : 
    (index==248) ? 32'h4017657d : 
    (index==249) ? 32'h40177fbb : 
    (index==250) ? 32'h401799fe : 
    (index==251) ? 32'h4017b446 : 
    (index==252) ? 32'h4017ce92 : 
    (index==253) ? 32'h4017e8e2 : 
    (index==254) ? 32'h40180338 : 
    (index==255) ? 32'h40181d91 : 
    (index==256) ? 32'h401837f0 : 
    (index==257) ? 32'h40185253 : 
    (index==258) ? 32'h40186cba : 
    (index==259) ? 32'h40188726 : 
    (index==260) ? 32'h4018a197 : 
    (index==261) ? 32'h4018bc0c : 
    (index==262) ? 32'h4018d686 : 
    (index==263) ? 32'h4018f104 : 
    (index==264) ? 32'h40190b87 : 
    (index==265) ? 32'h4019260f : 
    (index==266) ? 32'h4019409b : 
    (index==267) ? 32'h40195b2c : 
    (index==268) ? 32'h401975c1 : 
    (index==269) ? 32'h4019905b : 
    (index==270) ? 32'h4019aafa : 
    (index==271) ? 32'h4019c59d : 
    (index==272) ? 32'h4019e045 : 
    (index==273) ? 32'h4019faf2 : 
    (index==274) ? 32'h401a15a3 : 
    (index==275) ? 32'h401a3058 : 
    (index==276) ? 32'h401a4b13 : 
    (index==277) ? 32'h401a65d2 : 
    (index==278) ? 32'h401a8095 : 
    (index==279) ? 32'h401a9b5e : 
    (index==280) ? 32'h401ab62a : 
    (index==281) ? 32'h401ad0fc : 
    (index==282) ? 32'h401aebd2 : 
    (index==283) ? 32'h401b06ad : 
    (index==284) ? 32'h401b218d : 
    (index==285) ? 32'h401b3c71 : 
    (index==286) ? 32'h401b575a : 
    (index==287) ? 32'h401b7247 : 
    (index==288) ? 32'h401b8d39 : 
    (index==289) ? 32'h401ba830 : 
    (index==290) ? 32'h401bc32c : 
    (index==291) ? 32'h401bde2c : 
    (index==292) ? 32'h401bf931 : 
    (index==293) ? 32'h401c143a : 
    (index==294) ? 32'h401c2f48 : 
    (index==295) ? 32'h401c4a5b : 
    (index==296) ? 32'h401c6573 : 
    (index==297) ? 32'h401c808f : 
    (index==298) ? 32'h401c9bb0 : 
    (index==299) ? 32'h401cb6d6 : 
    (index==300) ? 32'h401cd200 : 
    (index==301) ? 32'h401ced2f : 
    (index==302) ? 32'h401d0863 : 
    (index==303) ? 32'h401d239c : 
    (index==304) ? 32'h401d3ed9 : 
    (index==305) ? 32'h401d5a1b : 
    (index==306) ? 32'h401d7562 : 
    (index==307) ? 32'h401d90ad : 
    (index==308) ? 32'h401dabfd : 
    (index==309) ? 32'h401dc752 : 
    (index==310) ? 32'h401de2ac : 
    (index==311) ? 32'h401dfe0a : 
    (index==312) ? 32'h401e196e : 
    (index==313) ? 32'h401e34d5 : 
    (index==314) ? 32'h401e5042 : 
    (index==315) ? 32'h401e6bb4 : 
    (index==316) ? 32'h401e872a : 
    (index==317) ? 32'h401ea2a5 : 
    (index==318) ? 32'h401ebe24 : 
    (index==319) ? 32'h401ed9a9 : 
    (index==320) ? 32'h401ef532 : 
    (index==321) ? 32'h401f10c0 : 
    (index==322) ? 32'h401f2c53 : 
    (index==323) ? 32'h401f47ea : 
    (index==324) ? 32'h401f6386 : 
    (index==325) ? 32'h401f7f28 : 
    (index==326) ? 32'h401f9acd : 
    (index==327) ? 32'h401fb678 : 
    (index==328) ? 32'h401fd228 : 
    (index==329) ? 32'h401feddc : 
    (index==330) ? 32'h40200995 : 
    (index==331) ? 32'h40202553 : 
    (index==332) ? 32'h40204116 : 
    (index==333) ? 32'h40205cdd : 
    (index==334) ? 32'h402078a9 : 
    (index==335) ? 32'h4020947b : 
    (index==336) ? 32'h4020b051 : 
    (index==337) ? 32'h4020cc2b : 
    (index==338) ? 32'h4020e80b : 
    (index==339) ? 32'h402103ef : 
    (index==340) ? 32'h40211fd9 : 
    (index==341) ? 32'h40213bc7 : 
    (index==342) ? 32'h402157ba : 
    (index==343) ? 32'h402173b2 : 
    (index==344) ? 32'h40218fae : 
    (index==345) ? 32'h4021abb0 : 
    (index==346) ? 32'h4021c7b6 : 
    (index==347) ? 32'h4021e3c1 : 
    (index==348) ? 32'h4021ffd1 : 
    (index==349) ? 32'h40221be6 : 
    (index==350) ? 32'h40223800 : 
    (index==351) ? 32'h4022541f : 
    (index==352) ? 32'h40227043 : 
    (index==353) ? 32'h40228c6b : 
    (index==354) ? 32'h4022a898 : 
    (index==355) ? 32'h4022c4ca : 
    (index==356) ? 32'h4022e102 : 
    (index==357) ? 32'h4022fd3e : 
    (index==358) ? 32'h4023197e : 
    (index==359) ? 32'h402335c4 : 
    (index==360) ? 32'h4023520f : 
    (index==361) ? 32'h40236e5e : 
    (index==362) ? 32'h40238ab3 : 
    (index==363) ? 32'h4023a70c : 
    (index==364) ? 32'h4023c36b : 
    (index==365) ? 32'h4023dfce : 
    (index==366) ? 32'h4023fc36 : 
    (index==367) ? 32'h402418a3 : 
    (index==368) ? 32'h40243515 : 
    (index==369) ? 32'h4024518c : 
    (index==370) ? 32'h40246e08 : 
    (index==371) ? 32'h40248a89 : 
    (index==372) ? 32'h4024a70f : 
    (index==373) ? 32'h4024c399 : 
    (index==374) ? 32'h4024e029 : 
    (index==375) ? 32'h4024fcbd : 
    (index==376) ? 32'h40251957 : 
    (index==377) ? 32'h402535f6 : 
    (index==378) ? 32'h40255299 : 
    (index==379) ? 32'h40256f41 : 
    (index==380) ? 32'h40258bef : 
    (index==381) ? 32'h4025a8a1 : 
    (index==382) ? 32'h4025c559 : 
    (index==383) ? 32'h4025e215 : 
    (index==384) ? 32'h4025fed6 : 
    (index==385) ? 32'h40261b9c : 
    (index==386) ? 32'h40263868 : 
    (index==387) ? 32'h40265538 : 
    (index==388) ? 32'h4026720d : 
    (index==389) ? 32'h40268ee8 : 
    (index==390) ? 32'h4026abc7 : 
    (index==391) ? 32'h4026c8ab : 
    (index==392) ? 32'h4026e594 : 
    (index==393) ? 32'h40270283 : 
    (index==394) ? 32'h40271f76 : 
    (index==395) ? 32'h40273c6e : 
    (index==396) ? 32'h4027596c : 
    (index==397) ? 32'h4027766e : 
    (index==398) ? 32'h40279375 : 
    (index==399) ? 32'h4027b082 : 
    (index==400) ? 32'h4027cd93 : 
    (index==401) ? 32'h4027eaaa : 
    (index==402) ? 32'h402807c5 : 
    (index==403) ? 32'h402824e6 : 
    (index==404) ? 32'h4028420b : 
    (index==405) ? 32'h40285f36 : 
    (index==406) ? 32'h40287c66 : 
    (index==407) ? 32'h4028999b : 
    (index==408) ? 32'h4028b6d5 : 
    (index==409) ? 32'h4028d414 : 
    (index==410) ? 32'h4028f158 : 
    (index==411) ? 32'h40290ea1 : 
    (index==412) ? 32'h40292bef : 
    (index==413) ? 32'h40294942 : 
    (index==414) ? 32'h4029669a : 
    (index==415) ? 32'h402983f8 : 
    (index==416) ? 32'h4029a15a : 
    (index==417) ? 32'h4029bec2 : 
    (index==418) ? 32'h4029dc2e : 
    (index==419) ? 32'h4029f9a0 : 
    (index==420) ? 32'h402a1717 : 
    (index==421) ? 32'h402a3493 : 
    (index==422) ? 32'h402a5214 : 
    (index==423) ? 32'h402a6f9a : 
    (index==424) ? 32'h402a8d26 : 
    (index==425) ? 32'h402aaab6 : 
    (index==426) ? 32'h402ac84c : 
    (index==427) ? 32'h402ae5e7 : 
    (index==428) ? 32'h402b0386 : 
    (index==429) ? 32'h402b212b : 
    (index==430) ? 32'h402b3ed6 : 
    (index==431) ? 32'h402b5c85 : 
    (index==432) ? 32'h402b7a39 : 
    (index==433) ? 32'h402b97f3 : 
    (index==434) ? 32'h402bb5b1 : 
    (index==435) ? 32'h402bd375 : 
    (index==436) ? 32'h402bf13e : 
    (index==437) ? 32'h402c0f0d : 
    (index==438) ? 32'h402c2ce0 : 
    (index==439) ? 32'h402c4ab8 : 
    (index==440) ? 32'h402c6896 : 
    (index==441) ? 32'h402c8679 : 
    (index==442) ? 32'h402ca461 : 
    (index==443) ? 32'h402cc24e : 
    (index==444) ? 32'h402ce041 : 
    (index==445) ? 32'h402cfe38 : 
    (index==446) ? 32'h402d1c35 : 
    (index==447) ? 32'h402d3a37 : 
    (index==448) ? 32'h402d583e : 
    (index==449) ? 32'h402d764b : 
    (index==450) ? 32'h402d945c : 
    (index==451) ? 32'h402db273 : 
    (index==452) ? 32'h402dd08f : 
    (index==453) ? 32'h402deeb1 : 
    (index==454) ? 32'h402e0cd7 : 
    (index==455) ? 32'h402e2b03 : 
    (index==456) ? 32'h402e4934 : 
    (index==457) ? 32'h402e676a : 
    (index==458) ? 32'h402e85a5 : 
    (index==459) ? 32'h402ea3e6 : 
    (index==460) ? 32'h402ec22c : 
    (index==461) ? 32'h402ee077 : 
    (index==462) ? 32'h402efec8 : 
    (index==463) ? 32'h402f1d1d : 
    (index==464) ? 32'h402f3b78 : 
    (index==465) ? 32'h402f59d8 : 
    (index==466) ? 32'h402f783e : 
    (index==467) ? 32'h402f96a9 : 
    (index==468) ? 32'h402fb519 : 
    (index==469) ? 32'h402fd38e : 
    (index==470) ? 32'h402ff208 : 
    (index==471) ? 32'h40301088 : 
    (index==472) ? 32'h40302f0d : 
    (index==473) ? 32'h40304d98 : 
    (index==474) ? 32'h40306c27 : 
    (index==475) ? 32'h40308abc : 
    (index==476) ? 32'h4030a957 : 
    (index==477) ? 32'h4030c7f6 : 
    (index==478) ? 32'h4030e69b : 
    (index==479) ? 32'h40310545 : 
    (index==480) ? 32'h403123f5 : 
    (index==481) ? 32'h403142aa : 
    (index==482) ? 32'h40316164 : 
    (index==483) ? 32'h40318024 : 
    (index==484) ? 32'h40319ee8 : 
    (index==485) ? 32'h4031bdb3 : 
    (index==486) ? 32'h4031dc82 : 
    (index==487) ? 32'h4031fb57 : 
    (index==488) ? 32'h40321a31 : 
    (index==489) ? 32'h40323911 : 
    (index==490) ? 32'h403257f6 : 
    (index==491) ? 32'h403276e0 : 
    (index==492) ? 32'h403295cf : 
    (index==493) ? 32'h4032b4c4 : 
    (index==494) ? 32'h4032d3bf : 
    (index==495) ? 32'h4032f2be : 
    (index==496) ? 32'h403311c4 : 
    (index==497) ? 32'h403330ce : 
    (index==498) ? 32'h40334fde : 
    (index==499) ? 32'h40336ef3 : 
    (index==500) ? 32'h40338e0e : 
    (index==501) ? 32'h4033ad2e : 
    (index==502) ? 32'h4033cc53 : 
    (index==503) ? 32'h4033eb7e : 
    (index==504) ? 32'h40340aae : 
    (index==505) ? 32'h403429e4 : 
    (index==506) ? 32'h4034491f : 
    (index==507) ? 32'h4034685f : 
    (index==508) ? 32'h403487a5 : 
    (index==509) ? 32'h4034a6f0 : 
    (index==510) ? 32'h4034c641 : 
    (index==511) ? 32'h4034e597 : 
    (index==512) ? 32'h403504f3 : 
    (index==513) ? 32'h40352454 : 
    (index==514) ? 32'h403543ba : 
    (index==515) ? 32'h40356326 : 
    (index==516) ? 32'h40358297 : 
    (index==517) ? 32'h4035a20e : 
    (index==518) ? 32'h4035c18a : 
    (index==519) ? 32'h4035e10c : 
    (index==520) ? 32'h40360093 : 
    (index==521) ? 32'h40362020 : 
    (index==522) ? 32'h40363fb2 : 
    (index==523) ? 32'h40365f49 : 
    (index==524) ? 32'h40367ee6 : 
    (index==525) ? 32'h40369e89 : 
    (index==526) ? 32'h4036be31 : 
    (index==527) ? 32'h4036ddde : 
    (index==528) ? 32'h4036fd91 : 
    (index==529) ? 32'h40371d4a : 
    (index==530) ? 32'h40373d08 : 
    (index==531) ? 32'h40375ccb : 
    (index==532) ? 32'h40377c94 : 
    (index==533) ? 32'h40379c63 : 
    (index==534) ? 32'h4037bc37 : 
    (index==535) ? 32'h4037dc10 : 
    (index==536) ? 32'h4037fbef : 
    (index==537) ? 32'h40381bd4 : 
    (index==538) ? 32'h40383bbe : 
    (index==539) ? 32'h40385bae : 
    (index==540) ? 32'h40387ba3 : 
    (index==541) ? 32'h40389b9d : 
    (index==542) ? 32'h4038bb9e : 
    (index==543) ? 32'h4038dba3 : 
    (index==544) ? 32'h4038fbaf : 
    (index==545) ? 32'h40391bc0 : 
    (index==546) ? 32'h40393bd6 : 
    (index==547) ? 32'h40395bf2 : 
    (index==548) ? 32'h40397c14 : 
    (index==549) ? 32'h40399c3b : 
    (index==550) ? 32'h4039bc68 : 
    (index==551) ? 32'h4039dc9a : 
    (index==552) ? 32'h4039fcd2 : 
    (index==553) ? 32'h403a1d0f : 
    (index==554) ? 32'h403a3d52 : 
    (index==555) ? 32'h403a5d9b : 
    (index==556) ? 32'h403a7de9 : 
    (index==557) ? 32'h403a9e3d : 
    (index==558) ? 32'h403abe96 : 
    (index==559) ? 32'h403adef6 : 
    (index==560) ? 32'h403aff5a : 
    (index==561) ? 32'h403b1fc4 : 
    (index==562) ? 32'h403b4034 : 
    (index==563) ? 32'h403b60aa : 
    (index==564) ? 32'h403b8125 : 
    (index==565) ? 32'h403ba1a6 : 
    (index==566) ? 32'h403bc22c : 
    (index==567) ? 32'h403be2b8 : 
    (index==568) ? 32'h403c034a : 
    (index==569) ? 32'h403c23e1 : 
    (index==570) ? 32'h403c447e : 
    (index==571) ? 32'h403c6521 : 
    (index==572) ? 32'h403c85c9 : 
    (index==573) ? 32'h403ca677 : 
    (index==574) ? 32'h403cc72b : 
    (index==575) ? 32'h403ce7e4 : 
    (index==576) ? 32'h403d08a3 : 
    (index==577) ? 32'h403d2968 : 
    (index==578) ? 32'h403d4a32 : 
    (index==579) ? 32'h403d6b02 : 
    (index==580) ? 32'h403d8bd8 : 
    (index==581) ? 32'h403dacb3 : 
    (index==582) ? 32'h403dcd94 : 
    (index==583) ? 32'h403dee7b : 
    (index==584) ? 32'h403e0f68 : 
    (index==585) ? 32'h403e305a : 
    (index==586) ? 32'h403e5152 : 
    (index==587) ? 32'h403e724f : 
    (index==588) ? 32'h403e9353 : 
    (index==589) ? 32'h403eb45c : 
    (index==590) ? 32'h403ed56a : 
    (index==591) ? 32'h403ef67f : 
    (index==592) ? 32'h403f1799 : 
    (index==593) ? 32'h403f38b9 : 
    (index==594) ? 32'h403f59df : 
    (index==595) ? 32'h403f7b0a : 
    (index==596) ? 32'h403f9c3c : 
    (index==597) ? 32'h403fbd73 : 
    (index==598) ? 32'h403fdeaf : 
    (index==599) ? 32'h403ffff2 : 
    (index==600) ? 32'h4040213a : 
    (index==601) ? 32'h40404288 : 
    (index==602) ? 32'h404063dc : 
    (index==603) ? 32'h40408536 : 
    (index==604) ? 32'h4040a695 : 
    (index==605) ? 32'h4040c7fa : 
    (index==606) ? 32'h4040e965 : 
    (index==607) ? 32'h40410ad6 : 
    (index==608) ? 32'h40412c4c : 
    (index==609) ? 32'h40414dc9 : 
    (index==610) ? 32'h40416f4b : 
    (index==611) ? 32'h404190d3 : 
    (index==612) ? 32'h4041b260 : 
    (index==613) ? 32'h4041d3f4 : 
    (index==614) ? 32'h4041f58d : 
    (index==615) ? 32'h4042172d : 
    (index==616) ? 32'h404238d2 : 
    (index==617) ? 32'h40425a7d : 
    (index==618) ? 32'h40427c2d : 
    (index==619) ? 32'h40429de4 : 
    (index==620) ? 32'h4042bfa0 : 
    (index==621) ? 32'h4042e162 : 
    (index==622) ? 32'h4043032b : 
    (index==623) ? 32'h404324f9 : 
    (index==624) ? 32'h404346cc : 
    (index==625) ? 32'h404368a6 : 
    (index==626) ? 32'h40438a86 : 
    (index==627) ? 32'h4043ac6b : 
    (index==628) ? 32'h4043ce56 : 
    (index==629) ? 32'h4043f047 : 
    (index==630) ? 32'h4044123f : 
    (index==631) ? 32'h4044343b : 
    (index==632) ? 32'h4044563e : 
    (index==633) ? 32'h40447847 : 
    (index==634) ? 32'h40449a56 : 
    (index==635) ? 32'h4044bc6a : 
    (index==636) ? 32'h4044de85 : 
    (index==637) ? 32'h404500a5 : 
    (index==638) ? 32'h404522cb : 
    (index==639) ? 32'h404544f7 : 
    (index==640) ? 32'h4045672a : 
    (index==641) ? 32'h40458962 : 
    (index==642) ? 32'h4045aba0 : 
    (index==643) ? 32'h4045cde3 : 
    (index==644) ? 32'h4045f02d : 
    (index==645) ? 32'h4046127d : 
    (index==646) ? 32'h404634d3 : 
    (index==647) ? 32'h4046572f : 
    (index==648) ? 32'h40467990 : 
    (index==649) ? 32'h40469bf8 : 
    (index==650) ? 32'h4046be65 : 
    (index==651) ? 32'h4046e0d9 : 
    (index==652) ? 32'h40470352 : 
    (index==653) ? 32'h404725d2 : 
    (index==654) ? 32'h40474857 : 
    (index==655) ? 32'h40476ae3 : 
    (index==656) ? 32'h40478d74 : 
    (index==657) ? 32'h4047b00c : 
    (index==658) ? 32'h4047d2a9 : 
    (index==659) ? 32'h4047f54d : 
    (index==660) ? 32'h404817f6 : 
    (index==661) ? 32'h40483aa5 : 
    (index==662) ? 32'h40485d5b : 
    (index==663) ? 32'h40488016 : 
    (index==664) ? 32'h4048a2d8 : 
    (index==665) ? 32'h4048c59f : 
    (index==666) ? 32'h4048e86d : 
    (index==667) ? 32'h40490b40 : 
    (index==668) ? 32'h40492e1a : 
    (index==669) ? 32'h404950fa : 
    (index==670) ? 32'h404973df : 
    (index==671) ? 32'h404996cb : 
    (index==672) ? 32'h4049b9bd : 
    (index==673) ? 32'h4049dcb5 : 
    (index==674) ? 32'h4049ffb3 : 
    (index==675) ? 32'h404a22b7 : 
    (index==676) ? 32'h404a45c1 : 
    (index==677) ? 32'h404a68d1 : 
    (index==678) ? 32'h404a8be7 : 
    (index==679) ? 32'h404aaf03 : 
    (index==680) ? 32'h404ad226 : 
    (index==681) ? 32'h404af54e : 
    (index==682) ? 32'h404b187d : 
    (index==683) ? 32'h404b3bb2 : 
    (index==684) ? 32'h404b5eec : 
    (index==685) ? 32'h404b822d : 
    (index==686) ? 32'h404ba574 : 
    (index==687) ? 32'h404bc8c1 : 
    (index==688) ? 32'h404bec14 : 
    (index==689) ? 32'h404c0f6e : 
    (index==690) ? 32'h404c32cd : 
    (index==691) ? 32'h404c5633 : 
    (index==692) ? 32'h404c799f : 
    (index==693) ? 32'h404c9d11 : 
    (index==694) ? 32'h404cc089 : 
    (index==695) ? 32'h404ce407 : 
    (index==696) ? 32'h404d078b : 
    (index==697) ? 32'h404d2b16 : 
    (index==698) ? 32'h404d4ea6 : 
    (index==699) ? 32'h404d723d : 
    (index==700) ? 32'h404d95da : 
    (index==701) ? 32'h404db97d : 
    (index==702) ? 32'h404ddd26 : 
    (index==703) ? 32'h404e00d6 : 
    (index==704) ? 32'h404e248c : 
    (index==705) ? 32'h404e4847 : 
    (index==706) ? 32'h404e6c0a : 
    (index==707) ? 32'h404e8fd2 : 
    (index==708) ? 32'h404eb3a0 : 
    (index==709) ? 32'h404ed775 : 
    (index==710) ? 32'h404efb50 : 
    (index==711) ? 32'h404f1f31 : 
    (index==712) ? 32'h404f4318 : 
    (index==713) ? 32'h404f6706 : 
    (index==714) ? 32'h404f8afa : 
    (index==715) ? 32'h404faef4 : 
    (index==716) ? 32'h404fd2f4 : 
    (index==717) ? 32'h404ff6fa : 
    (index==718) ? 32'h40501b07 : 
    (index==719) ? 32'h40503f1a : 
    (index==720) ? 32'h40506333 : 
    (index==721) ? 32'h40508753 : 
    (index==722) ? 32'h4050ab79 : 
    (index==723) ? 32'h4050cfa5 : 
    (index==724) ? 32'h4050f3d7 : 
    (index==725) ? 32'h4051180f : 
    (index==726) ? 32'h40513c4e : 
    (index==727) ? 32'h40516093 : 
    (index==728) ? 32'h405184df : 
    (index==729) ? 32'h4051a931 : 
    (index==730) ? 32'h4051cd89 : 
    (index==731) ? 32'h4051f1e7 : 
    (index==732) ? 32'h4052164c : 
    (index==733) ? 32'h40523ab6 : 
    (index==734) ? 32'h40525f28 : 
    (index==735) ? 32'h4052839f : 
    (index==736) ? 32'h4052a81d : 
    (index==737) ? 32'h4052cca1 : 
    (index==738) ? 32'h4052f12c : 
    (index==739) ? 32'h405315bd : 
    (index==740) ? 32'h40533a54 : 
    (index==741) ? 32'h40535ef1 : 
    (index==742) ? 32'h40538395 : 
    (index==743) ? 32'h4053a840 : 
    (index==744) ? 32'h4053ccf0 : 
    (index==745) ? 32'h4053f1a7 : 
    (index==746) ? 32'h40541664 : 
    (index==747) ? 32'h40543b28 : 
    (index==748) ? 32'h40545ff2 : 
    (index==749) ? 32'h405484c3 : 
    (index==750) ? 32'h4054a999 : 
    (index==751) ? 32'h4054ce77 : 
    (index==752) ? 32'h4054f35a : 
    (index==753) ? 32'h40551844 : 
    (index==754) ? 32'h40553d35 : 
    (index==755) ? 32'h4055622b : 
    (index==756) ? 32'h40558729 : 
    (index==757) ? 32'h4055ac2c : 
    (index==758) ? 32'h4055d136 : 
    (index==759) ? 32'h4055f647 : 
    (index==760) ? 32'h40561b5d : 
    (index==761) ? 32'h4056407b : 
    (index==762) ? 32'h4056659f : 
    (index==763) ? 32'h40568ac9 : 
    (index==764) ? 32'h4056aff9 : 
    (index==765) ? 32'h4056d530 : 
    (index==766) ? 32'h4056fa6e : 
    (index==767) ? 32'h40571fb2 : 
    (index==768) ? 32'h405744fc : 
    (index==769) ? 32'h40576a4d : 
    (index==770) ? 32'h40578fa5 : 
    (index==771) ? 32'h4057b502 : 
    (index==772) ? 32'h4057da67 : 
    (index==773) ? 32'h4057ffd1 : 
    (index==774) ? 32'h40582543 : 
    (index==775) ? 32'h40584abb : 
    (index==776) ? 32'h40587039 : 
    (index==777) ? 32'h405895be : 
    (index==778) ? 32'h4058bb49 : 
    (index==779) ? 32'h4058e0db : 
    (index==780) ? 32'h40590673 : 
    (index==781) ? 32'h40592c12 : 
    (index==782) ? 32'h405951b7 : 
    (index==783) ? 32'h40597763 : 
    (index==784) ? 32'h40599d15 : 
    (index==785) ? 32'h4059c2ce : 
    (index==786) ? 32'h4059e88e : 
    (index==787) ? 32'h405a0e54 : 
    (index==788) ? 32'h405a3420 : 
    (index==789) ? 32'h405a59f3 : 
    (index==790) ? 32'h405a7fcd : 
    (index==791) ? 32'h405aa5ad : 
    (index==792) ? 32'h405acb94 : 
    (index==793) ? 32'h405af181 : 
    (index==794) ? 32'h405b1775 : 
    (index==795) ? 32'h405b3d70 : 
    (index==796) ? 32'h405b6371 : 
    (index==797) ? 32'h405b8978 : 
    (index==798) ? 32'h405baf87 : 
    (index==799) ? 32'h405bd59c : 
    (index==800) ? 32'h405bfbb7 : 
    (index==801) ? 32'h405c21d9 : 
    (index==802) ? 32'h405c4802 : 
    (index==803) ? 32'h405c6e31 : 
    (index==804) ? 32'h405c9467 : 
    (index==805) ? 32'h405cbaa4 : 
    (index==806) ? 32'h405ce0e7 : 
    (index==807) ? 32'h405d0731 : 
    (index==808) ? 32'h405d2d81 : 
    (index==809) ? 32'h405d53d8 : 
    (index==810) ? 32'h405d7a36 : 
    (index==811) ? 32'h405da09a : 
    (index==812) ? 32'h405dc705 : 
    (index==813) ? 32'h405ded77 : 
    (index==814) ? 32'h405e13ef : 
    (index==815) ? 32'h405e3a6e : 
    (index==816) ? 32'h405e60f4 : 
    (index==817) ? 32'h405e8780 : 
    (index==818) ? 32'h405eae13 : 
    (index==819) ? 32'h405ed4ad : 
    (index==820) ? 32'h405efb4e : 
    (index==821) ? 32'h405f21f5 : 
    (index==822) ? 32'h405f48a3 : 
    (index==823) ? 32'h405f6f57 : 
    (index==824) ? 32'h405f9612 : 
    (index==825) ? 32'h405fbcd4 : 
    (index==826) ? 32'h405fe39d : 
    (index==827) ? 32'h40600a6c : 
    (index==828) ? 32'h40603143 : 
    (index==829) ? 32'h4060581f : 
    (index==830) ? 32'h40607f03 : 
    (index==831) ? 32'h4060a5ed : 
    (index==832) ? 32'h4060ccde : 
    (index==833) ? 32'h4060f3d6 : 
    (index==834) ? 32'h40611ad5 : 
    (index==835) ? 32'h406141da : 
    (index==836) ? 32'h406168e6 : 
    (index==837) ? 32'h40618ff9 : 
    (index==838) ? 32'h4061b713 : 
    (index==839) ? 32'h4061de33 : 
    (index==840) ? 32'h4062055a : 
    (index==841) ? 32'h40622c89 : 
    (index==842) ? 32'h406253bd : 
    (index==843) ? 32'h40627af9 : 
    (index==844) ? 32'h4062a23b : 
    (index==845) ? 32'h4062c984 : 
    (index==846) ? 32'h4062f0d4 : 
    (index==847) ? 32'h4063182b : 
    (index==848) ? 32'h40633f89 : 
    (index==849) ? 32'h406366ed : 
    (index==850) ? 32'h40638e59 : 
    (index==851) ? 32'h4063b5cb : 
    (index==852) ? 32'h4063dd44 : 
    (index==853) ? 32'h406404c4 : 
    (index==854) ? 32'h40642c4a : 
    (index==855) ? 32'h406453d8 : 
    (index==856) ? 32'h40647b6c : 
    (index==857) ? 32'h4064a307 : 
    (index==858) ? 32'h4064caa9 : 
    (index==859) ? 32'h4064f252 : 
    (index==860) ? 32'h40651a02 : 
    (index==861) ? 32'h406541b9 : 
    (index==862) ? 32'h40656977 : 
    (index==863) ? 32'h4065913b : 
    (index==864) ? 32'h4065b906 : 
    (index==865) ? 32'h4065e0d9 : 
    (index==866) ? 32'h406608b2 : 
    (index==867) ? 32'h40663092 : 
    (index==868) ? 32'h40665879 : 
    (index==869) ? 32'h40668067 : 
    (index==870) ? 32'h4066a85c : 
    (index==871) ? 32'h4066d057 : 
    (index==872) ? 32'h4066f85a : 
    (index==873) ? 32'h40672064 : 
    (index==874) ? 32'h40674874 : 
    (index==875) ? 32'h4067708c : 
    (index==876) ? 32'h406798aa : 
    (index==877) ? 32'h4067c0d0 : 
    (index==878) ? 32'h4067e8fc : 
    (index==879) ? 32'h40681130 : 
    (index==880) ? 32'h4068396a : 
    (index==881) ? 32'h406861ab : 
    (index==882) ? 32'h406889f3 : 
    (index==883) ? 32'h4068b243 : 
    (index==884) ? 32'h4068da99 : 
    (index==885) ? 32'h406902f6 : 
    (index==886) ? 32'h40692b5a : 
    (index==887) ? 32'h406953c6 : 
    (index==888) ? 32'h40697c38 : 
    (index==889) ? 32'h4069a4b1 : 
    (index==890) ? 32'h4069cd31 : 
    (index==891) ? 32'h4069f5b9 : 
    (index==892) ? 32'h406a1e47 : 
    (index==893) ? 32'h406a46dc : 
    (index==894) ? 32'h406a6f79 : 
    (index==895) ? 32'h406a981c : 
    (index==896) ? 32'h406ac0c6 : 
    (index==897) ? 32'h406ae978 : 
    (index==898) ? 32'h406b1230 : 
    (index==899) ? 32'h406b3af0 : 
    (index==900) ? 32'h406b63b7 : 
    (index==901) ? 32'h406b8c85 : 
    (index==902) ? 32'h406bb559 : 
    (index==903) ? 32'h406bde35 : 
    (index==904) ? 32'h406c0718 : 
    (index==905) ? 32'h406c3002 : 
    (index==906) ? 32'h406c58f3 : 
    (index==907) ? 32'h406c81ec : 
    (index==908) ? 32'h406caaeb : 
    (index==909) ? 32'h406cd3f2 : 
    (index==910) ? 32'h406cfcff : 
    (index==911) ? 32'h406d2614 : 
    (index==912) ? 32'h406d4f30 : 
    (index==913) ? 32'h406d7853 : 
    (index==914) ? 32'h406da17d : 
    (index==915) ? 32'h406dcaae : 
    (index==916) ? 32'h406df3e6 : 
    (index==917) ? 32'h406e1d26 : 
    (index==918) ? 32'h406e466c : 
    (index==919) ? 32'h406e6fba : 
    (index==920) ? 32'h406e990f : 
    (index==921) ? 32'h406ec26b : 
    (index==922) ? 32'h406eebcf : 
    (index==923) ? 32'h406f1539 : 
    (index==924) ? 32'h406f3eab : 
    (index==925) ? 32'h406f6823 : 
    (index==926) ? 32'h406f91a3 : 
    (index==927) ? 32'h406fbb2b : 
    (index==928) ? 32'h406fe4b9 : 
    (index==929) ? 32'h40700e4f : 
    (index==930) ? 32'h407037ec : 
    (index==931) ? 32'h40706190 : 
    (index==932) ? 32'h40708b3b : 
    (index==933) ? 32'h4070b4ed : 
    (index==934) ? 32'h4070dea7 : 
    (index==935) ? 32'h40710868 : 
    (index==936) ? 32'h40713230 : 
    (index==937) ? 32'h40715c00 : 
    (index==938) ? 32'h407185d6 : 
    (index==939) ? 32'h4071afb4 : 
    (index==940) ? 32'h4071d999 : 
    (index==941) ? 32'h40720386 : 
    (index==942) ? 32'h40722d79 : 
    (index==943) ? 32'h40725774 : 
    (index==944) ? 32'h40728177 : 
    (index==945) ? 32'h4072ab80 : 
    (index==946) ? 32'h4072d591 : 
    (index==947) ? 32'h4072ffa9 : 
    (index==948) ? 32'h407329c9 : 
    (index==949) ? 32'h407353ef : 
    (index==950) ? 32'h40737e1d : 
    (index==951) ? 32'h4073a853 : 
    (index==952) ? 32'h4073d28f : 
    (index==953) ? 32'h4073fcd3 : 
    (index==954) ? 32'h4074271f : 
    (index==955) ? 32'h40745171 : 
    (index==956) ? 32'h40747bcb : 
    (index==957) ? 32'h4074a62d : 
    (index==958) ? 32'h4074d095 : 
    (index==959) ? 32'h4074fb05 : 
    (index==960) ? 32'h4075257d : 
    (index==961) ? 32'h40754ffb : 
    (index==962) ? 32'h40757a81 : 
    (index==963) ? 32'h4075a50f : 
    (index==964) ? 32'h4075cfa4 : 
    (index==965) ? 32'h4075fa40 : 
    (index==966) ? 32'h407624e4 : 
    (index==967) ? 32'h40764f8f : 
    (index==968) ? 32'h40767a41 : 
    (index==969) ? 32'h4076a4fb : 
    (index==970) ? 32'h4076cfbc : 
    (index==971) ? 32'h4076fa85 : 
    (index==972) ? 32'h40772555 : 
    (index==973) ? 32'h4077502c : 
    (index==974) ? 32'h40777b0b : 
    (index==975) ? 32'h4077a5f1 : 
    (index==976) ? 32'h4077d0df : 
    (index==977) ? 32'h4077fbd4 : 
    (index==978) ? 32'h407826d1 : 
    (index==979) ? 32'h407851d5 : 
    (index==980) ? 32'h40787ce0 : 
    (index==981) ? 32'h4078a7f3 : 
    (index==982) ? 32'h4078d30e : 
    (index==983) ? 32'h4078fe30 : 
    (index==984) ? 32'h40792959 : 
    (index==985) ? 32'h4079548a : 
    (index==986) ? 32'h40797fc3 : 
    (index==987) ? 32'h4079ab02 : 
    (index==988) ? 32'h4079d64a : 
    (index==989) ? 32'h407a0199 : 
    (index==990) ? 32'h407a2cef : 
    (index==991) ? 32'h407a584d : 
    (index==992) ? 32'h407a83b2 : 
    (index==993) ? 32'h407aaf1f : 
    (index==994) ? 32'h407ada94 : 
    (index==995) ? 32'h407b0610 : 
    (index==996) ? 32'h407b3193 : 
    (index==997) ? 32'h407b5d1e : 
    (index==998) ? 32'h407b88b1 : 
    (index==999) ? 32'h407bb44b : 
    (index==1000) ? 32'h407bdfed : 
    (index==1001) ? 32'h407c0b96 : 
    (index==1002) ? 32'h407c3747 : 
    (index==1003) ? 32'h407c6300 : 
    (index==1004) ? 32'h407c8ec0 : 
    (index==1005) ? 32'h407cba87 : 
    (index==1006) ? 32'h407ce656 : 
    (index==1007) ? 32'h407d122d : 
    (index==1008) ? 32'h407d3e0c : 
    (index==1009) ? 32'h407d69f2 : 
    (index==1010) ? 32'h407d95df : 
    (index==1011) ? 32'h407dc1d4 : 
    (index==1012) ? 32'h407dedd1 : 
    (index==1013) ? 32'h407e19d6 : 
    (index==1014) ? 32'h407e45e2 : 
    (index==1015) ? 32'h407e71f5 : 
    (index==1016) ? 32'h407e9e11 : 
    (index==1017) ? 32'h407eca34 : 
    (index==1018) ? 32'h407ef65f : 
    (index==1019) ? 32'h407f2291 : 
    (index==1020) ? 32'h407f4ecb : 
    (index==1021) ? 32'h407f7b0c : 
    (index==1022) ? 32'h407fa756 : 
    (index==1023) ? 32'h407fd3a7 : 
    0;
endmodule
