module Flt_sqrt_u40_5(
    input [39:0] ain
    ,input  clk
    ,input  en
    ,output  [19:0] out
    ,input  rst_n
    ,input  vldin
    ,output   vldout
);
wire  vld20;
wire [39:0] datain20;
wire [39:0] Y20;
wire [39:0] YY20;
wire [39:0] Decra19;
wire [39:0] Decrb19;
wire [39:0] Decr19;
wire [39:0] YY19_1;
wire [39:0] Base19;
wire  smaller19;
wire [39:0] YY19;
wire [19:0] Y19;
wire [39:0] datain19;
wire  vld19;
wire [39:0] Decra18;
wire [39:0] Decrb18;
wire [39:0] Decr18;
wire [39:0] YY18_1;
wire [39:0] Base18;
wire  smaller18;
wire [39:0] YY18;
wire [19:0] Y18;
wire [39:0] datain18;
wire  vld18;
wire [39:0] Decra17;
wire [39:0] Decrb17;
wire [39:0] Decr17;
wire [39:0] YY17_1;
wire [39:0] Base17;
wire  smaller17;
wire [39:0] YY17;
wire [19:0] Y17;
wire [39:0] datain17;
wire  vld17;
wire [39:0] Decra16;
wire [39:0] Decrb16;
wire [39:0] Decr16;
wire [39:0] YY16_1;
wire [39:0] Base16;
wire  smaller16;
wire [39:0] YY16;
wire [19:0] Y16;
wire [39:0] datain16;
wire  vld16;
wire [39:0] Decra15;
wire [39:0] Decrb15;
wire [39:0] Decr15;
wire [39:0] YY15_1;
wire [39:0] Base15;
wire  smaller15;
wire [39:0] pre_YY15;
wire [19:0] pre_Y15;
wire [39:0] YY15;
wire [39:0] Y15;
wire [39:0] datain15;
wire  vld15;
wire [39:0] Decra14;
wire [39:0] Decrb14;
wire [39:0] Decr14;
wire [39:0] YY14_1;
wire [39:0] Base14;
wire  smaller14;
wire [39:0] YY14;
wire [19:0] Y14;
wire [39:0] datain14;
wire  vld14;
wire [39:0] Decra13;
wire [39:0] Decrb13;
wire [39:0] Decr13;
wire [39:0] YY13_1;
wire [39:0] Base13;
wire  smaller13;
wire [39:0] YY13;
wire [19:0] Y13;
wire [39:0] datain13;
wire  vld13;
wire [39:0] Decra12;
wire [39:0] Decrb12;
wire [39:0] Decr12;
wire [39:0] YY12_1;
wire [39:0] Base12;
wire  smaller12;
wire [39:0] YY12;
wire [19:0] Y12;
wire [39:0] datain12;
wire  vld12;
wire [39:0] Decra11;
wire [39:0] Decrb11;
wire [39:0] Decr11;
wire [39:0] YY11_1;
wire [39:0] Base11;
wire  smaller11;
wire [39:0] YY11;
wire [19:0] Y11;
wire [39:0] datain11;
wire  vld11;
wire [39:0] Decra10;
wire [39:0] Decrb10;
wire [39:0] Decr10;
wire [39:0] YY10_1;
wire [39:0] Base10;
wire  smaller10;
wire [39:0] pre_YY10;
wire [19:0] pre_Y10;
wire [39:0] YY10;
wire [39:0] Y10;
wire [39:0] datain10;
wire  vld10;
wire [39:0] Decra9;
wire [39:0] Decrb9;
wire [39:0] Decr9;
wire [39:0] YY9_1;
wire [39:0] Base9;
wire  smaller9;
wire [39:0] YY9;
wire [19:0] Y9;
wire [39:0] datain9;
wire  vld9;
wire [39:0] Decra8;
wire [39:0] Decrb8;
wire [39:0] Decr8;
wire [39:0] YY8_1;
wire [39:0] Base8;
wire  smaller8;
wire [39:0] YY8;
wire [19:0] Y8;
wire [39:0] datain8;
wire  vld8;
wire [39:0] Decra7;
wire [39:0] Decrb7;
wire [39:0] Decr7;
wire [39:0] YY7_1;
wire [39:0] Base7;
wire  smaller7;
wire [39:0] YY7;
wire [19:0] Y7;
wire [39:0] datain7;
wire  vld7;
wire [39:0] Decra6;
wire [39:0] Decrb6;
wire [39:0] Decr6;
wire [39:0] YY6_1;
wire [39:0] Base6;
wire  smaller6;
wire [39:0] YY6;
wire [19:0] Y6;
wire [39:0] datain6;
wire  vld6;
wire [39:0] Decra5;
wire [39:0] Decrb5;
wire [39:0] Decr5;
wire [39:0] YY5_1;
wire [39:0] Base5;
wire  smaller5;
wire [39:0] pre_YY5;
wire [19:0] pre_Y5;
wire [39:0] YY5;
wire [39:0] Y5;
wire [39:0] datain5;
wire  vld5;
wire [39:0] Decra4;
wire [39:0] Decrb4;
wire [39:0] Decr4;
wire [39:0] YY4_1;
wire [39:0] Base4;
wire  smaller4;
wire [39:0] YY4;
wire [19:0] Y4;
wire [39:0] datain4;
wire  vld4;
wire [39:0] Decra3;
wire [39:0] Decrb3;
wire [39:0] Decr3;
wire [39:0] YY3_1;
wire [39:0] Base3;
wire  smaller3;
wire [39:0] YY3;
wire [19:0] Y3;
wire [39:0] datain3;
wire  vld3;
wire [39:0] Decra2;
wire [39:0] Decrb2;
wire [39:0] Decr2;
wire [39:0] YY2_1;
wire [39:0] Base2;
wire  smaller2;
wire [39:0] YY2;
wire [19:0] Y2;
wire [39:0] datain2;
wire  vld2;
wire [39:0] Decra1;
wire [39:0] Decrb1;
wire [39:0] Decr1;
wire [39:0] YY1_1;
wire [39:0] Base1;
wire  smaller1;
wire [39:0] YY1;
wire [19:0] Y1;
wire [39:0] datain1;
wire  vld1;
wire [39:0] Decra0;
wire [39:0] Decrb0;
wire [39:0] Decr0;
wire [39:0] YY0_1;
wire [39:0] Base0;
wire  smaller0;
wire [39:0] YY0;
wire [19:0] Y0;
wire [39:0] datain0;
wire  vld0;
wire [39:0] Flt_Y20;
wire [39:0] Flt_YY20;
wire [39:0] Flt_Decra19;
wire [39:0] Flt_Decrb19;
wire [39:0] Flt_Decr19;
wire [39:0] Flt_YY19_1;
wire [39:0] Flt_Base19;
wire  Flt_smaller19;
wire [39:0] Flt_YY19;
wire [19:0] Flt_Y19;
wire [39:0] Flt_datain19;
wire  Flt_vld19;
wire [39:0] Flt_Decra18;
wire [39:0] Flt_Decrb18;
wire [39:0] Flt_Decr18;
wire [39:0] Flt_YY18_1;
wire [39:0] Flt_Base18;
wire  Flt_smaller18;
wire [39:0] Flt_YY18;
wire [19:0] Flt_Y18;
wire [39:0] Flt_datain18;
wire  Flt_vld18;
wire [39:0] Flt_Decra17;
wire [39:0] Flt_Decrb17;
wire [39:0] Flt_Decr17;
wire [39:0] Flt_YY17_1;
wire [39:0] Flt_Base17;
wire  Flt_smaller17;
wire [39:0] Flt_YY17;
wire [19:0] Flt_Y17;
wire [39:0] Flt_datain17;
wire  Flt_vld17;
wire [39:0] Flt_Decra16;
wire [39:0] Flt_Decrb16;
wire [39:0] Flt_Decr16;
wire [39:0] Flt_YY16_1;
wire [39:0] Flt_Base16;
wire  Flt_smaller16;
wire [39:0] Flt_YY16;
wire [19:0] Flt_Y16;
wire [39:0] Flt_datain16;
wire  Flt_vld16;
wire [39:0] Flt_Decra15;
wire [39:0] Flt_Decrb15;
wire [39:0] Flt_Decr15;
wire [39:0] Flt_YY15_1;
wire [39:0] Flt_Base15;
wire  Flt_smaller15;
wire [39:0] Flt_pre_YY15;
wire [19:0] Flt_pre_Y15;
wire [39:0] Flt_Decra14;
wire [39:0] Flt_Decrb14;
wire [39:0] Flt_Decr14;
wire [39:0] Flt_YY14_1;
wire [39:0] Flt_Base14;
wire  Flt_smaller14;
wire [39:0] Flt_YY14;
wire [19:0] Flt_Y14;
wire [39:0] Flt_datain14;
wire  Flt_vld14;
wire [39:0] Flt_Decra13;
wire [39:0] Flt_Decrb13;
wire [39:0] Flt_Decr13;
wire [39:0] Flt_YY13_1;
wire [39:0] Flt_Base13;
wire  Flt_smaller13;
wire [39:0] Flt_YY13;
wire [19:0] Flt_Y13;
wire [39:0] Flt_datain13;
wire  Flt_vld13;
wire [39:0] Flt_Decra12;
wire [39:0] Flt_Decrb12;
wire [39:0] Flt_Decr12;
wire [39:0] Flt_YY12_1;
wire [39:0] Flt_Base12;
wire  Flt_smaller12;
wire [39:0] Flt_YY12;
wire [19:0] Flt_Y12;
wire [39:0] Flt_datain12;
wire  Flt_vld12;
wire [39:0] Flt_Decra11;
wire [39:0] Flt_Decrb11;
wire [39:0] Flt_Decr11;
wire [39:0] Flt_YY11_1;
wire [39:0] Flt_Base11;
wire  Flt_smaller11;
wire [39:0] Flt_YY11;
wire [19:0] Flt_Y11;
wire [39:0] Flt_datain11;
wire  Flt_vld11;
wire [39:0] Flt_Decra10;
wire [39:0] Flt_Decrb10;
wire [39:0] Flt_Decr10;
wire [39:0] Flt_YY10_1;
wire [39:0] Flt_Base10;
wire  Flt_smaller10;
wire [39:0] Flt_pre_YY10;
wire [19:0] Flt_pre_Y10;
wire [39:0] Flt_Decra9;
wire [39:0] Flt_Decrb9;
wire [39:0] Flt_Decr9;
wire [39:0] Flt_YY9_1;
wire [39:0] Flt_Base9;
wire  Flt_smaller9;
wire [39:0] Flt_YY9;
wire [19:0] Flt_Y9;
wire [39:0] Flt_datain9;
wire  Flt_vld9;
wire [39:0] Flt_Decra8;
wire [39:0] Flt_Decrb8;
wire [39:0] Flt_Decr8;
wire [39:0] Flt_YY8_1;
wire [39:0] Flt_Base8;
wire  Flt_smaller8;
wire [39:0] Flt_YY8;
wire [19:0] Flt_Y8;
wire [39:0] Flt_datain8;
wire  Flt_vld8;
wire [39:0] Flt_Decra7;
wire [39:0] Flt_Decrb7;
wire [39:0] Flt_Decr7;
wire [39:0] Flt_YY7_1;
wire [39:0] Flt_Base7;
wire  Flt_smaller7;
wire [39:0] Flt_YY7;
wire [19:0] Flt_Y7;
wire [39:0] Flt_datain7;
wire  Flt_vld7;
wire [39:0] Flt_Decra6;
wire [39:0] Flt_Decrb6;
wire [39:0] Flt_Decr6;
wire [39:0] Flt_YY6_1;
wire [39:0] Flt_Base6;
wire  Flt_smaller6;
wire [39:0] Flt_YY6;
wire [19:0] Flt_Y6;
wire [39:0] Flt_datain6;
wire  Flt_vld6;
wire [39:0] Flt_Decra5;
wire [39:0] Flt_Decrb5;
wire [39:0] Flt_Decr5;
wire [39:0] Flt_YY5_1;
wire [39:0] Flt_Base5;
wire  Flt_smaller5;
wire [39:0] Flt_pre_YY5;
wire [19:0] Flt_pre_Y5;
wire [39:0] Flt_Decra4;
wire [39:0] Flt_Decrb4;
wire [39:0] Flt_Decr4;
wire [39:0] Flt_YY4_1;
wire [39:0] Flt_Base4;
wire  Flt_smaller4;
wire [39:0] Flt_YY4;
wire [19:0] Flt_Y4;
wire [39:0] Flt_datain4;
wire  Flt_vld4;
wire [39:0] Flt_Decra3;
wire [39:0] Flt_Decrb3;
wire [39:0] Flt_Decr3;
wire [39:0] Flt_YY3_1;
wire [39:0] Flt_Base3;
wire  Flt_smaller3;
wire [39:0] Flt_YY3;
wire [19:0] Flt_Y3;
wire [39:0] Flt_datain3;
wire  Flt_vld3;
wire [39:0] Flt_Decra2;
wire [39:0] Flt_Decrb2;
wire [39:0] Flt_Decr2;
wire [39:0] Flt_YY2_1;
wire [39:0] Flt_Base2;
wire  Flt_smaller2;
wire [39:0] Flt_YY2;
wire [19:0] Flt_Y2;
wire [39:0] Flt_datain2;
wire  Flt_vld2;
wire [39:0] Flt_Decra1;
wire [39:0] Flt_Decrb1;
wire [39:0] Flt_Decr1;
wire [39:0] Flt_YY1_1;
wire [39:0] Flt_Base1;
wire  Flt_smaller1;
wire [39:0] Flt_YY1;
wire [19:0] Flt_Y1;
wire [39:0] Flt_datain1;
wire  Flt_vld1;
wire [39:0] Flt_Decra0;
wire [39:0] Flt_Decrb0;
wire [39:0] Flt_Decr0;
wire [39:0] Flt_YY0_1;
wire [39:0] Flt_Base0;
wire  Flt_smaller0;
wire [39:0] Flt_YY0;
wire [19:0] Flt_Y0;
wire [39:0] Flt_datain0;
wire  Flt_vld0;
reg  Flt_vld20;
reg [39:0] Flt_datain20;
reg [39:0] Flt_YY15;
reg [39:0] Flt_Y15;
reg [39:0] Flt_datain15;
reg  Flt_vld15;
reg [39:0] Flt_YY10;
reg [39:0] Flt_Y10;
reg [39:0] Flt_datain10;
reg  Flt_vld10;
reg [39:0] Flt_YY5;
reg [39:0] Flt_Y5;
reg [39:0] Flt_datain5;
reg  Flt_vld5;
reg [19:0] Flt_out;
reg  Flt_vldout;
assign   Flt_Y20 = 0;
assign   Flt_YY20 = 0;
assign   Flt_Decra19 = 40'b1 << 38;
assign   Flt_Decrb19 = Y20 << 20;
assign   Flt_Decr19 = Decra19 + Decrb19;
assign   Flt_YY19_1 = YY20 + Decr19;
assign   Flt_Base19 = 40'b1 << 19;
assign   Flt_smaller19 = YY19_1 <= datain20;
assign   Flt_YY19 = smaller19 ? YY19_1 : YY20;
assign   Flt_Y19 = smaller19 ? (Y20 + Base19) : Y20;
assign   Flt_datain19 = datain20;
assign   Flt_vld19 = vld20;
assign   Flt_Decra18 = 40'b1 << 36;
assign   Flt_Decrb18 = Y19 << 19;
assign   Flt_Decr18 = Decra18 + Decrb18;
assign   Flt_YY18_1 = YY19 + Decr18;
assign   Flt_Base18 = 40'b1 << 18;
assign   Flt_smaller18 = YY18_1 <= datain19;
assign   Flt_YY18 = smaller18 ? YY18_1 : YY19;
assign   Flt_Y18 = smaller18 ? (Y19 + Base18) : Y19;
assign   Flt_datain18 = datain19;
assign   Flt_vld18 = vld19;
assign   Flt_Decra17 = 40'b1 << 34;
assign   Flt_Decrb17 = Y18 << 18;
assign   Flt_Decr17 = Decra17 + Decrb17;
assign   Flt_YY17_1 = YY18 + Decr17;
assign   Flt_Base17 = 40'b1 << 17;
assign   Flt_smaller17 = YY17_1 <= datain18;
assign   Flt_YY17 = smaller17 ? YY17_1 : YY18;
assign   Flt_Y17 = smaller17 ? (Y18 + Base17) : Y18;
assign   Flt_datain17 = datain18;
assign   Flt_vld17 = vld18;
assign   Flt_Decra16 = 40'b1 << 32;
assign   Flt_Decrb16 = Y17 << 17;
assign   Flt_Decr16 = Decra16 + Decrb16;
assign   Flt_YY16_1 = YY17 + Decr16;
assign   Flt_Base16 = 40'b1 << 16;
assign   Flt_smaller16 = YY16_1 <= datain17;
assign   Flt_YY16 = smaller16 ? YY16_1 : YY17;
assign   Flt_Y16 = smaller16 ? (Y17 + Base16) : Y17;
assign   Flt_datain16 = datain17;
assign   Flt_vld16 = vld17;
assign   Flt_Decra15 = 40'b1 << 30;
assign   Flt_Decrb15 = Y16 << 16;
assign   Flt_Decr15 = Decra15 + Decrb15;
assign   Flt_YY15_1 = YY16 + Decr15;
assign   Flt_Base15 = 40'b1 << 15;
assign   Flt_smaller15 = YY15_1 <= datain16;
assign   Flt_pre_YY15 = smaller15 ? YY15_1 : YY16;
assign   Flt_pre_Y15 = smaller15 ? (Y16 + Base15) : Y16;
assign   Flt_Decra14 = 40'b1 << 28;
assign   Flt_Decrb14 = Y15 << 15;
assign   Flt_Decr14 = Decra14 + Decrb14;
assign   Flt_YY14_1 = YY15 + Decr14;
assign   Flt_Base14 = 40'b1 << 14;
assign   Flt_smaller14 = YY14_1 <= datain15;
assign   Flt_YY14 = smaller14 ? YY14_1 : YY15;
assign   Flt_Y14 = smaller14 ? (Y15 + Base14) : Y15;
assign   Flt_datain14 = datain15;
assign   Flt_vld14 = vld15;
assign   Flt_Decra13 = 40'b1 << 26;
assign   Flt_Decrb13 = Y14 << 14;
assign   Flt_Decr13 = Decra13 + Decrb13;
assign   Flt_YY13_1 = YY14 + Decr13;
assign   Flt_Base13 = 40'b1 << 13;
assign   Flt_smaller13 = YY13_1 <= datain14;
assign   Flt_YY13 = smaller13 ? YY13_1 : YY14;
assign   Flt_Y13 = smaller13 ? (Y14 + Base13) : Y14;
assign   Flt_datain13 = datain14;
assign   Flt_vld13 = vld14;
assign   Flt_Decra12 = 40'b1 << 24;
assign   Flt_Decrb12 = Y13 << 13;
assign   Flt_Decr12 = Decra12 + Decrb12;
assign   Flt_YY12_1 = YY13 + Decr12;
assign   Flt_Base12 = 40'b1 << 12;
assign   Flt_smaller12 = YY12_1 <= datain13;
assign   Flt_YY12 = smaller12 ? YY12_1 : YY13;
assign   Flt_Y12 = smaller12 ? (Y13 + Base12) : Y13;
assign   Flt_datain12 = datain13;
assign   Flt_vld12 = vld13;
assign   Flt_Decra11 = 40'b1 << 22;
assign   Flt_Decrb11 = Y12 << 12;
assign   Flt_Decr11 = Decra11 + Decrb11;
assign   Flt_YY11_1 = YY12 + Decr11;
assign   Flt_Base11 = 40'b1 << 11;
assign   Flt_smaller11 = YY11_1 <= datain12;
assign   Flt_YY11 = smaller11 ? YY11_1 : YY12;
assign   Flt_Y11 = smaller11 ? (Y12 + Base11) : Y12;
assign   Flt_datain11 = datain12;
assign   Flt_vld11 = vld12;
assign   Flt_Decra10 = 40'b1 << 20;
assign   Flt_Decrb10 = Y11 << 11;
assign   Flt_Decr10 = Decra10 + Decrb10;
assign   Flt_YY10_1 = YY11 + Decr10;
assign   Flt_Base10 = 40'b1 << 10;
assign   Flt_smaller10 = YY10_1 <= datain11;
assign   Flt_pre_YY10 = smaller10 ? YY10_1 : YY11;
assign   Flt_pre_Y10 = smaller10 ? (Y11 + Base10) : Y11;
assign   Flt_Decra9 = 40'b1 << 18;
assign   Flt_Decrb9 = Y10 << 10;
assign   Flt_Decr9 = Decra9 + Decrb9;
assign   Flt_YY9_1 = YY10 + Decr9;
assign   Flt_Base9 = 40'b1 << 9;
assign   Flt_smaller9 = YY9_1 <= datain10;
assign   Flt_YY9 = smaller9 ? YY9_1 : YY10;
assign   Flt_Y9 = smaller9 ? (Y10 + Base9) : Y10;
assign   Flt_datain9 = datain10;
assign   Flt_vld9 = vld10;
assign   Flt_Decra8 = 40'b1 << 16;
assign   Flt_Decrb8 = Y9 << 9;
assign   Flt_Decr8 = Decra8 + Decrb8;
assign   Flt_YY8_1 = YY9 + Decr8;
assign   Flt_Base8 = 40'b1 << 8;
assign   Flt_smaller8 = YY8_1 <= datain9;
assign   Flt_YY8 = smaller8 ? YY8_1 : YY9;
assign   Flt_Y8 = smaller8 ? (Y9 + Base8) : Y9;
assign   Flt_datain8 = datain9;
assign   Flt_vld8 = vld9;
assign   Flt_Decra7 = 40'b1 << 14;
assign   Flt_Decrb7 = Y8 << 8;
assign   Flt_Decr7 = Decra7 + Decrb7;
assign   Flt_YY7_1 = YY8 + Decr7;
assign   Flt_Base7 = 40'b1 << 7;
assign   Flt_smaller7 = YY7_1 <= datain8;
assign   Flt_YY7 = smaller7 ? YY7_1 : YY8;
assign   Flt_Y7 = smaller7 ? (Y8 + Base7) : Y8;
assign   Flt_datain7 = datain8;
assign   Flt_vld7 = vld8;
assign   Flt_Decra6 = 40'b1 << 12;
assign   Flt_Decrb6 = Y7 << 7;
assign   Flt_Decr6 = Decra6 + Decrb6;
assign   Flt_YY6_1 = YY7 + Decr6;
assign   Flt_Base6 = 40'b1 << 6;
assign   Flt_smaller6 = YY6_1 <= datain7;
assign   Flt_YY6 = smaller6 ? YY6_1 : YY7;
assign   Flt_Y6 = smaller6 ? (Y7 + Base6) : Y7;
assign   Flt_datain6 = datain7;
assign   Flt_vld6 = vld7;
assign   Flt_Decra5 = 40'b1 << 10;
assign   Flt_Decrb5 = Y6 << 6;
assign   Flt_Decr5 = Decra5 + Decrb5;
assign   Flt_YY5_1 = YY6 + Decr5;
assign   Flt_Base5 = 40'b1 << 5;
assign   Flt_smaller5 = YY5_1 <= datain6;
assign   Flt_pre_YY5 = smaller5 ? YY5_1 : YY6;
assign   Flt_pre_Y5 = smaller5 ? (Y6 + Base5) : Y6;
assign   Flt_Decra4 = 40'b1 << 8;
assign   Flt_Decrb4 = Y5 << 5;
assign   Flt_Decr4 = Decra4 + Decrb4;
assign   Flt_YY4_1 = YY5 + Decr4;
assign   Flt_Base4 = 40'b1 << 4;
assign   Flt_smaller4 = YY4_1 <= datain5;
assign   Flt_YY4 = smaller4 ? YY4_1 : YY5;
assign   Flt_Y4 = smaller4 ? (Y5 + Base4) : Y5;
assign   Flt_datain4 = datain5;
assign   Flt_vld4 = vld5;
assign   Flt_Decra3 = 40'b1 << 6;
assign   Flt_Decrb3 = Y4 << 4;
assign   Flt_Decr3 = Decra3 + Decrb3;
assign   Flt_YY3_1 = YY4 + Decr3;
assign   Flt_Base3 = 40'b1 << 3;
assign   Flt_smaller3 = YY3_1 <= datain4;
assign   Flt_YY3 = smaller3 ? YY3_1 : YY4;
assign   Flt_Y3 = smaller3 ? (Y4 + Base3) : Y4;
assign   Flt_datain3 = datain4;
assign   Flt_vld3 = vld4;
assign   Flt_Decra2 = 40'b1 << 4;
assign   Flt_Decrb2 = Y3 << 3;
assign   Flt_Decr2 = Decra2 + Decrb2;
assign   Flt_YY2_1 = YY3 + Decr2;
assign   Flt_Base2 = 40'b1 << 2;
assign   Flt_smaller2 = YY2_1 <= datain3;
assign   Flt_YY2 = smaller2 ? YY2_1 : YY3;
assign   Flt_Y2 = smaller2 ? (Y3 + Base2) : Y3;
assign   Flt_datain2 = datain3;
assign   Flt_vld2 = vld3;
assign   Flt_Decra1 = 40'b1 << 2;
assign   Flt_Decrb1 = Y2 << 2;
assign   Flt_Decr1 = Decra1 + Decrb1;
assign   Flt_YY1_1 = YY2 + Decr1;
assign   Flt_Base1 = 40'b1 << 1;
assign   Flt_smaller1 = YY1_1 <= datain2;
assign   Flt_YY1 = smaller1 ? YY1_1 : YY2;
assign   Flt_Y1 = smaller1 ? (Y2 + Base1) : Y2;
assign   Flt_datain1 = datain2;
assign   Flt_vld1 = vld2;
assign   Flt_Decra0 = 40'b1 << 0;
assign   Flt_Decrb0 = Y1 << 1;
assign   Flt_Decr0 = Decra0 + Decrb0;
assign   Flt_YY0_1 = YY1 + Decr0;
assign   Flt_Base0 = 40'b1 << 0;
assign   Flt_smaller0 = YY0_1 <= datain1;
assign   Flt_YY0 = smaller0 ? YY0_1 : YY1;
assign   Flt_Y0 = smaller0 ? (Y1 + Base0) : Y1;
assign   Flt_datain0 = datain1;
assign   Flt_vld0 = vld1;
faultifizer #(.WID(40)) faultify_Y20 (.inx(Flt_Y20), .outx(Y20));
faultifizer #(.WID(40)) faultify_YY20 (.inx(Flt_YY20), .outx(YY20));
faultifizer #(.WID(40)) faultify_Decra19 (.inx(Flt_Decra19), .outx(Decra19));
faultifizer #(.WID(40)) faultify_Decrb19 (.inx(Flt_Decrb19), .outx(Decrb19));
faultifizer #(.WID(40)) faultify_Decr19 (.inx(Flt_Decr19), .outx(Decr19));
faultifizer #(.WID(40)) faultify_YY19_1 (.inx(Flt_YY19_1), .outx(YY19_1));
faultifizer #(.WID(40)) faultify_Base19 (.inx(Flt_Base19), .outx(Base19));
faultifizer #(.WID(1)) faultify_smaller19 (.inx(Flt_smaller19), .outx(smaller19));
faultifizer #(.WID(40)) faultify_YY19 (.inx(Flt_YY19), .outx(YY19));
faultifizer #(.WID(20)) faultify_Y19 (.inx(Flt_Y19), .outx(Y19));
faultifizer #(.WID(40)) faultify_datain19 (.inx(Flt_datain19), .outx(datain19));
faultifizer #(.WID(1)) faultify_vld19 (.inx(Flt_vld19), .outx(vld19));
faultifizer #(.WID(40)) faultify_Decra18 (.inx(Flt_Decra18), .outx(Decra18));
faultifizer #(.WID(40)) faultify_Decrb18 (.inx(Flt_Decrb18), .outx(Decrb18));
faultifizer #(.WID(40)) faultify_Decr18 (.inx(Flt_Decr18), .outx(Decr18));
faultifizer #(.WID(40)) faultify_YY18_1 (.inx(Flt_YY18_1), .outx(YY18_1));
faultifizer #(.WID(40)) faultify_Base18 (.inx(Flt_Base18), .outx(Base18));
faultifizer #(.WID(1)) faultify_smaller18 (.inx(Flt_smaller18), .outx(smaller18));
faultifizer #(.WID(40)) faultify_YY18 (.inx(Flt_YY18), .outx(YY18));
faultifizer #(.WID(20)) faultify_Y18 (.inx(Flt_Y18), .outx(Y18));
faultifizer #(.WID(40)) faultify_datain18 (.inx(Flt_datain18), .outx(datain18));
faultifizer #(.WID(1)) faultify_vld18 (.inx(Flt_vld18), .outx(vld18));
faultifizer #(.WID(40)) faultify_Decra17 (.inx(Flt_Decra17), .outx(Decra17));
faultifizer #(.WID(40)) faultify_Decrb17 (.inx(Flt_Decrb17), .outx(Decrb17));
faultifizer #(.WID(40)) faultify_Decr17 (.inx(Flt_Decr17), .outx(Decr17));
faultifizer #(.WID(40)) faultify_YY17_1 (.inx(Flt_YY17_1), .outx(YY17_1));
faultifizer #(.WID(40)) faultify_Base17 (.inx(Flt_Base17), .outx(Base17));
faultifizer #(.WID(1)) faultify_smaller17 (.inx(Flt_smaller17), .outx(smaller17));
faultifizer #(.WID(40)) faultify_YY17 (.inx(Flt_YY17), .outx(YY17));
faultifizer #(.WID(20)) faultify_Y17 (.inx(Flt_Y17), .outx(Y17));
faultifizer #(.WID(40)) faultify_datain17 (.inx(Flt_datain17), .outx(datain17));
faultifizer #(.WID(1)) faultify_vld17 (.inx(Flt_vld17), .outx(vld17));
faultifizer #(.WID(40)) faultify_Decra16 (.inx(Flt_Decra16), .outx(Decra16));
faultifizer #(.WID(40)) faultify_Decrb16 (.inx(Flt_Decrb16), .outx(Decrb16));
faultifizer #(.WID(40)) faultify_Decr16 (.inx(Flt_Decr16), .outx(Decr16));
faultifizer #(.WID(40)) faultify_YY16_1 (.inx(Flt_YY16_1), .outx(YY16_1));
faultifizer #(.WID(40)) faultify_Base16 (.inx(Flt_Base16), .outx(Base16));
faultifizer #(.WID(1)) faultify_smaller16 (.inx(Flt_smaller16), .outx(smaller16));
faultifizer #(.WID(40)) faultify_YY16 (.inx(Flt_YY16), .outx(YY16));
faultifizer #(.WID(20)) faultify_Y16 (.inx(Flt_Y16), .outx(Y16));
faultifizer #(.WID(40)) faultify_datain16 (.inx(Flt_datain16), .outx(datain16));
faultifizer #(.WID(1)) faultify_vld16 (.inx(Flt_vld16), .outx(vld16));
faultifizer #(.WID(40)) faultify_Decra15 (.inx(Flt_Decra15), .outx(Decra15));
faultifizer #(.WID(40)) faultify_Decrb15 (.inx(Flt_Decrb15), .outx(Decrb15));
faultifizer #(.WID(40)) faultify_Decr15 (.inx(Flt_Decr15), .outx(Decr15));
faultifizer #(.WID(40)) faultify_YY15_1 (.inx(Flt_YY15_1), .outx(YY15_1));
faultifizer #(.WID(40)) faultify_Base15 (.inx(Flt_Base15), .outx(Base15));
faultifizer #(.WID(1)) faultify_smaller15 (.inx(Flt_smaller15), .outx(smaller15));
faultifizer #(.WID(40)) faultify_pre_YY15 (.inx(Flt_pre_YY15), .outx(pre_YY15));
faultifizer #(.WID(20)) faultify_pre_Y15 (.inx(Flt_pre_Y15), .outx(pre_Y15));
faultifizer #(.WID(40)) faultify_Decra14 (.inx(Flt_Decra14), .outx(Decra14));
faultifizer #(.WID(40)) faultify_Decrb14 (.inx(Flt_Decrb14), .outx(Decrb14));
faultifizer #(.WID(40)) faultify_Decr14 (.inx(Flt_Decr14), .outx(Decr14));
faultifizer #(.WID(40)) faultify_YY14_1 (.inx(Flt_YY14_1), .outx(YY14_1));
faultifizer #(.WID(40)) faultify_Base14 (.inx(Flt_Base14), .outx(Base14));
faultifizer #(.WID(1)) faultify_smaller14 (.inx(Flt_smaller14), .outx(smaller14));
faultifizer #(.WID(40)) faultify_YY14 (.inx(Flt_YY14), .outx(YY14));
faultifizer #(.WID(20)) faultify_Y14 (.inx(Flt_Y14), .outx(Y14));
faultifizer #(.WID(40)) faultify_datain14 (.inx(Flt_datain14), .outx(datain14));
faultifizer #(.WID(1)) faultify_vld14 (.inx(Flt_vld14), .outx(vld14));
faultifizer #(.WID(40)) faultify_Decra13 (.inx(Flt_Decra13), .outx(Decra13));
faultifizer #(.WID(40)) faultify_Decrb13 (.inx(Flt_Decrb13), .outx(Decrb13));
faultifizer #(.WID(40)) faultify_Decr13 (.inx(Flt_Decr13), .outx(Decr13));
faultifizer #(.WID(40)) faultify_YY13_1 (.inx(Flt_YY13_1), .outx(YY13_1));
faultifizer #(.WID(40)) faultify_Base13 (.inx(Flt_Base13), .outx(Base13));
faultifizer #(.WID(1)) faultify_smaller13 (.inx(Flt_smaller13), .outx(smaller13));
faultifizer #(.WID(40)) faultify_YY13 (.inx(Flt_YY13), .outx(YY13));
faultifizer #(.WID(20)) faultify_Y13 (.inx(Flt_Y13), .outx(Y13));
faultifizer #(.WID(40)) faultify_datain13 (.inx(Flt_datain13), .outx(datain13));
faultifizer #(.WID(1)) faultify_vld13 (.inx(Flt_vld13), .outx(vld13));
faultifizer #(.WID(40)) faultify_Decra12 (.inx(Flt_Decra12), .outx(Decra12));
faultifizer #(.WID(40)) faultify_Decrb12 (.inx(Flt_Decrb12), .outx(Decrb12));
faultifizer #(.WID(40)) faultify_Decr12 (.inx(Flt_Decr12), .outx(Decr12));
faultifizer #(.WID(40)) faultify_YY12_1 (.inx(Flt_YY12_1), .outx(YY12_1));
faultifizer #(.WID(40)) faultify_Base12 (.inx(Flt_Base12), .outx(Base12));
faultifizer #(.WID(1)) faultify_smaller12 (.inx(Flt_smaller12), .outx(smaller12));
faultifizer #(.WID(40)) faultify_YY12 (.inx(Flt_YY12), .outx(YY12));
faultifizer #(.WID(20)) faultify_Y12 (.inx(Flt_Y12), .outx(Y12));
faultifizer #(.WID(40)) faultify_datain12 (.inx(Flt_datain12), .outx(datain12));
faultifizer #(.WID(1)) faultify_vld12 (.inx(Flt_vld12), .outx(vld12));
faultifizer #(.WID(40)) faultify_Decra11 (.inx(Flt_Decra11), .outx(Decra11));
faultifizer #(.WID(40)) faultify_Decrb11 (.inx(Flt_Decrb11), .outx(Decrb11));
faultifizer #(.WID(40)) faultify_Decr11 (.inx(Flt_Decr11), .outx(Decr11));
faultifizer #(.WID(40)) faultify_YY11_1 (.inx(Flt_YY11_1), .outx(YY11_1));
faultifizer #(.WID(40)) faultify_Base11 (.inx(Flt_Base11), .outx(Base11));
faultifizer #(.WID(1)) faultify_smaller11 (.inx(Flt_smaller11), .outx(smaller11));
faultifizer #(.WID(40)) faultify_YY11 (.inx(Flt_YY11), .outx(YY11));
faultifizer #(.WID(20)) faultify_Y11 (.inx(Flt_Y11), .outx(Y11));
faultifizer #(.WID(40)) faultify_datain11 (.inx(Flt_datain11), .outx(datain11));
faultifizer #(.WID(1)) faultify_vld11 (.inx(Flt_vld11), .outx(vld11));
faultifizer #(.WID(40)) faultify_Decra10 (.inx(Flt_Decra10), .outx(Decra10));
faultifizer #(.WID(40)) faultify_Decrb10 (.inx(Flt_Decrb10), .outx(Decrb10));
faultifizer #(.WID(40)) faultify_Decr10 (.inx(Flt_Decr10), .outx(Decr10));
faultifizer #(.WID(40)) faultify_YY10_1 (.inx(Flt_YY10_1), .outx(YY10_1));
faultifizer #(.WID(40)) faultify_Base10 (.inx(Flt_Base10), .outx(Base10));
faultifizer #(.WID(1)) faultify_smaller10 (.inx(Flt_smaller10), .outx(smaller10));
faultifizer #(.WID(40)) faultify_pre_YY10 (.inx(Flt_pre_YY10), .outx(pre_YY10));
faultifizer #(.WID(20)) faultify_pre_Y10 (.inx(Flt_pre_Y10), .outx(pre_Y10));
faultifizer #(.WID(40)) faultify_Decra9 (.inx(Flt_Decra9), .outx(Decra9));
faultifizer #(.WID(40)) faultify_Decrb9 (.inx(Flt_Decrb9), .outx(Decrb9));
faultifizer #(.WID(40)) faultify_Decr9 (.inx(Flt_Decr9), .outx(Decr9));
faultifizer #(.WID(40)) faultify_YY9_1 (.inx(Flt_YY9_1), .outx(YY9_1));
faultifizer #(.WID(40)) faultify_Base9 (.inx(Flt_Base9), .outx(Base9));
faultifizer #(.WID(1)) faultify_smaller9 (.inx(Flt_smaller9), .outx(smaller9));
faultifizer #(.WID(40)) faultify_YY9 (.inx(Flt_YY9), .outx(YY9));
faultifizer #(.WID(20)) faultify_Y9 (.inx(Flt_Y9), .outx(Y9));
faultifizer #(.WID(40)) faultify_datain9 (.inx(Flt_datain9), .outx(datain9));
faultifizer #(.WID(1)) faultify_vld9 (.inx(Flt_vld9), .outx(vld9));
faultifizer #(.WID(40)) faultify_Decra8 (.inx(Flt_Decra8), .outx(Decra8));
faultifizer #(.WID(40)) faultify_Decrb8 (.inx(Flt_Decrb8), .outx(Decrb8));
faultifizer #(.WID(40)) faultify_Decr8 (.inx(Flt_Decr8), .outx(Decr8));
faultifizer #(.WID(40)) faultify_YY8_1 (.inx(Flt_YY8_1), .outx(YY8_1));
faultifizer #(.WID(40)) faultify_Base8 (.inx(Flt_Base8), .outx(Base8));
faultifizer #(.WID(1)) faultify_smaller8 (.inx(Flt_smaller8), .outx(smaller8));
faultifizer #(.WID(40)) faultify_YY8 (.inx(Flt_YY8), .outx(YY8));
faultifizer #(.WID(20)) faultify_Y8 (.inx(Flt_Y8), .outx(Y8));
faultifizer #(.WID(40)) faultify_datain8 (.inx(Flt_datain8), .outx(datain8));
faultifizer #(.WID(1)) faultify_vld8 (.inx(Flt_vld8), .outx(vld8));
faultifizer #(.WID(40)) faultify_Decra7 (.inx(Flt_Decra7), .outx(Decra7));
faultifizer #(.WID(40)) faultify_Decrb7 (.inx(Flt_Decrb7), .outx(Decrb7));
faultifizer #(.WID(40)) faultify_Decr7 (.inx(Flt_Decr7), .outx(Decr7));
faultifizer #(.WID(40)) faultify_YY7_1 (.inx(Flt_YY7_1), .outx(YY7_1));
faultifizer #(.WID(40)) faultify_Base7 (.inx(Flt_Base7), .outx(Base7));
faultifizer #(.WID(1)) faultify_smaller7 (.inx(Flt_smaller7), .outx(smaller7));
faultifizer #(.WID(40)) faultify_YY7 (.inx(Flt_YY7), .outx(YY7));
faultifizer #(.WID(20)) faultify_Y7 (.inx(Flt_Y7), .outx(Y7));
faultifizer #(.WID(40)) faultify_datain7 (.inx(Flt_datain7), .outx(datain7));
faultifizer #(.WID(1)) faultify_vld7 (.inx(Flt_vld7), .outx(vld7));
faultifizer #(.WID(40)) faultify_Decra6 (.inx(Flt_Decra6), .outx(Decra6));
faultifizer #(.WID(40)) faultify_Decrb6 (.inx(Flt_Decrb6), .outx(Decrb6));
faultifizer #(.WID(40)) faultify_Decr6 (.inx(Flt_Decr6), .outx(Decr6));
faultifizer #(.WID(40)) faultify_YY6_1 (.inx(Flt_YY6_1), .outx(YY6_1));
faultifizer #(.WID(40)) faultify_Base6 (.inx(Flt_Base6), .outx(Base6));
faultifizer #(.WID(1)) faultify_smaller6 (.inx(Flt_smaller6), .outx(smaller6));
faultifizer #(.WID(40)) faultify_YY6 (.inx(Flt_YY6), .outx(YY6));
faultifizer #(.WID(20)) faultify_Y6 (.inx(Flt_Y6), .outx(Y6));
faultifizer #(.WID(40)) faultify_datain6 (.inx(Flt_datain6), .outx(datain6));
faultifizer #(.WID(1)) faultify_vld6 (.inx(Flt_vld6), .outx(vld6));
faultifizer #(.WID(40)) faultify_Decra5 (.inx(Flt_Decra5), .outx(Decra5));
faultifizer #(.WID(40)) faultify_Decrb5 (.inx(Flt_Decrb5), .outx(Decrb5));
faultifizer #(.WID(40)) faultify_Decr5 (.inx(Flt_Decr5), .outx(Decr5));
faultifizer #(.WID(40)) faultify_YY5_1 (.inx(Flt_YY5_1), .outx(YY5_1));
faultifizer #(.WID(40)) faultify_Base5 (.inx(Flt_Base5), .outx(Base5));
faultifizer #(.WID(1)) faultify_smaller5 (.inx(Flt_smaller5), .outx(smaller5));
faultifizer #(.WID(40)) faultify_pre_YY5 (.inx(Flt_pre_YY5), .outx(pre_YY5));
faultifizer #(.WID(20)) faultify_pre_Y5 (.inx(Flt_pre_Y5), .outx(pre_Y5));
faultifizer #(.WID(40)) faultify_Decra4 (.inx(Flt_Decra4), .outx(Decra4));
faultifizer #(.WID(40)) faultify_Decrb4 (.inx(Flt_Decrb4), .outx(Decrb4));
faultifizer #(.WID(40)) faultify_Decr4 (.inx(Flt_Decr4), .outx(Decr4));
faultifizer #(.WID(40)) faultify_YY4_1 (.inx(Flt_YY4_1), .outx(YY4_1));
faultifizer #(.WID(40)) faultify_Base4 (.inx(Flt_Base4), .outx(Base4));
faultifizer #(.WID(1)) faultify_smaller4 (.inx(Flt_smaller4), .outx(smaller4));
faultifizer #(.WID(40)) faultify_YY4 (.inx(Flt_YY4), .outx(YY4));
faultifizer #(.WID(20)) faultify_Y4 (.inx(Flt_Y4), .outx(Y4));
faultifizer #(.WID(40)) faultify_datain4 (.inx(Flt_datain4), .outx(datain4));
faultifizer #(.WID(1)) faultify_vld4 (.inx(Flt_vld4), .outx(vld4));
faultifizer #(.WID(40)) faultify_Decra3 (.inx(Flt_Decra3), .outx(Decra3));
faultifizer #(.WID(40)) faultify_Decrb3 (.inx(Flt_Decrb3), .outx(Decrb3));
faultifizer #(.WID(40)) faultify_Decr3 (.inx(Flt_Decr3), .outx(Decr3));
faultifizer #(.WID(40)) faultify_YY3_1 (.inx(Flt_YY3_1), .outx(YY3_1));
faultifizer #(.WID(40)) faultify_Base3 (.inx(Flt_Base3), .outx(Base3));
faultifizer #(.WID(1)) faultify_smaller3 (.inx(Flt_smaller3), .outx(smaller3));
faultifizer #(.WID(40)) faultify_YY3 (.inx(Flt_YY3), .outx(YY3));
faultifizer #(.WID(20)) faultify_Y3 (.inx(Flt_Y3), .outx(Y3));
faultifizer #(.WID(40)) faultify_datain3 (.inx(Flt_datain3), .outx(datain3));
faultifizer #(.WID(1)) faultify_vld3 (.inx(Flt_vld3), .outx(vld3));
faultifizer #(.WID(40)) faultify_Decra2 (.inx(Flt_Decra2), .outx(Decra2));
faultifizer #(.WID(40)) faultify_Decrb2 (.inx(Flt_Decrb2), .outx(Decrb2));
faultifizer #(.WID(40)) faultify_Decr2 (.inx(Flt_Decr2), .outx(Decr2));
faultifizer #(.WID(40)) faultify_YY2_1 (.inx(Flt_YY2_1), .outx(YY2_1));
faultifizer #(.WID(40)) faultify_Base2 (.inx(Flt_Base2), .outx(Base2));
faultifizer #(.WID(1)) faultify_smaller2 (.inx(Flt_smaller2), .outx(smaller2));
faultifizer #(.WID(40)) faultify_YY2 (.inx(Flt_YY2), .outx(YY2));
faultifizer #(.WID(20)) faultify_Y2 (.inx(Flt_Y2), .outx(Y2));
faultifizer #(.WID(40)) faultify_datain2 (.inx(Flt_datain2), .outx(datain2));
faultifizer #(.WID(1)) faultify_vld2 (.inx(Flt_vld2), .outx(vld2));
faultifizer #(.WID(40)) faultify_Decra1 (.inx(Flt_Decra1), .outx(Decra1));
faultifizer #(.WID(40)) faultify_Decrb1 (.inx(Flt_Decrb1), .outx(Decrb1));
faultifizer #(.WID(40)) faultify_Decr1 (.inx(Flt_Decr1), .outx(Decr1));
faultifizer #(.WID(40)) faultify_YY1_1 (.inx(Flt_YY1_1), .outx(YY1_1));
faultifizer #(.WID(40)) faultify_Base1 (.inx(Flt_Base1), .outx(Base1));
faultifizer #(.WID(1)) faultify_smaller1 (.inx(Flt_smaller1), .outx(smaller1));
faultifizer #(.WID(40)) faultify_YY1 (.inx(Flt_YY1), .outx(YY1));
faultifizer #(.WID(20)) faultify_Y1 (.inx(Flt_Y1), .outx(Y1));
faultifizer #(.WID(40)) faultify_datain1 (.inx(Flt_datain1), .outx(datain1));
faultifizer #(.WID(1)) faultify_vld1 (.inx(Flt_vld1), .outx(vld1));
faultifizer #(.WID(40)) faultify_Decra0 (.inx(Flt_Decra0), .outx(Decra0));
faultifizer #(.WID(40)) faultify_Decrb0 (.inx(Flt_Decrb0), .outx(Decrb0));
faultifizer #(.WID(40)) faultify_Decr0 (.inx(Flt_Decr0), .outx(Decr0));
faultifizer #(.WID(40)) faultify_YY0_1 (.inx(Flt_YY0_1), .outx(YY0_1));
faultifizer #(.WID(40)) faultify_Base0 (.inx(Flt_Base0), .outx(Base0));
faultifizer #(.WID(1)) faultify_smaller0 (.inx(Flt_smaller0), .outx(smaller0));
faultifizer #(.WID(40)) faultify_YY0 (.inx(Flt_YY0), .outx(YY0));
faultifizer #(.WID(20)) faultify_Y0 (.inx(Flt_Y0), .outx(Y0));
faultifizer #(.WID(40)) faultify_datain0 (.inx(Flt_datain0), .outx(datain0));
faultifizer #(.WID(1)) faultify_vld0 (.inx(Flt_vld0), .outx(vld0));
faultifizer #(.WID(1)) faultify_vld20 (.inx(Flt_vld20), .outx(vld20));
faultifizer #(.WID(40)) faultify_datain20 (.inx(Flt_datain20), .outx(datain20));
faultifizer #(.WID(40)) faultify_YY15 (.inx(Flt_YY15), .outx(YY15));
faultifizer #(.WID(40)) faultify_Y15 (.inx(Flt_Y15), .outx(Y15));
faultifizer #(.WID(40)) faultify_datain15 (.inx(Flt_datain15), .outx(datain15));
faultifizer #(.WID(1)) faultify_vld15 (.inx(Flt_vld15), .outx(vld15));
faultifizer #(.WID(40)) faultify_YY10 (.inx(Flt_YY10), .outx(YY10));
faultifizer #(.WID(40)) faultify_Y10 (.inx(Flt_Y10), .outx(Y10));
faultifizer #(.WID(40)) faultify_datain10 (.inx(Flt_datain10), .outx(datain10));
faultifizer #(.WID(1)) faultify_vld10 (.inx(Flt_vld10), .outx(vld10));
faultifizer #(.WID(40)) faultify_YY5 (.inx(Flt_YY5), .outx(YY5));
faultifizer #(.WID(40)) faultify_Y5 (.inx(Flt_Y5), .outx(Y5));
faultifizer #(.WID(40)) faultify_datain5 (.inx(Flt_datain5), .outx(datain5));
faultifizer #(.WID(1)) faultify_vld5 (.inx(Flt_vld5), .outx(vld5));
faultifizer #(.WID(20)) faultify_out (.inx(Flt_out), .outx(out));
faultifizer #(.WID(1)) faultify_vldout (.inx(Flt_vldout), .outx(vldout));
always @(posedge clk) begin
    if(en) begin
        Flt_vld20 <= vldin;
    end
end
always @(posedge clk) begin
    if(en) begin
        Flt_datain20 <= ain;
    end
end
always @(posedge clk) begin
    if(en) begin
        Flt_YY15 <= pre_YY15;
    end
end
always @(posedge clk) begin
    if(en) begin
        Flt_Y15 <= pre_Y15;
    end
end
always @(posedge clk) begin
    if(en) begin
        Flt_datain15 <= datain16;
    end
end
always @(posedge clk) begin
    if(en) begin
        Flt_vld15 <= vld16;
    end
end
always @(posedge clk) begin
    if(en) begin
        Flt_YY10 <= pre_YY10;
    end
end
always @(posedge clk) begin
    if(en) begin
        Flt_Y10 <= pre_Y10;
    end
end
always @(posedge clk) begin
    if(en) begin
        Flt_datain10 <= datain11;
    end
end
always @(posedge clk) begin
    if(en) begin
        Flt_vld10 <= vld11;
    end
end
always @(posedge clk) begin
    if(en) begin
        Flt_YY5 <= pre_YY5;
    end
end
always @(posedge clk) begin
    if(en) begin
        Flt_Y5 <= pre_Y5;
    end
end
always @(posedge clk) begin
    if(en) begin
        Flt_datain5 <= datain6;
    end
end
always @(posedge clk) begin
    if(en) begin
        Flt_vld5 <= vld6;
    end
end
always @(posedge clk) begin
    if(en) begin
        Flt_out <= Y0;
    end
end
always @(posedge clk) begin
    if(en) begin
        Flt_vldout <= vld0;
    end
end
endmodule

