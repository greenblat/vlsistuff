`timescale 1ns/1ps
module tb;
reg [31:0] cycles;   initial cycles=0;
reg [31:0] errors;   initial errors=0;
reg [31:0] wrongs;   initial wrongs=0;
reg [31:0] panics;   initial panics=0;
reg [31:0] corrects; initial corrects=0;
reg [31:0] marker;   initial marker=0;
reg [31:0] marker0;   initial marker0=0;
reg [31:0] marker1;   initial marker1=0;
reg [31:0] marker2;   initial marker2=0;
reg [31:0] marker3;   initial marker3=0;
reg [31:0] Index;   initial Index=0;


reg [2:0] mst0_awsize; initial mst0_awsize=3;
reg [2:0] mst1_awsize; initial mst1_awsize=3;
reg [2:0] mst2_awsize; initial mst2_awsize=3;
reg [2:0] mst3_awsize; initial mst3_awsize=3;

reg [2:0] mst0_arsize; initial mst0_arsize=3;
reg [2:0] mst1_arsize; initial mst1_arsize=3;
reg [2:0] mst2_arsize; initial mst2_arsize=3;
reg [2:0] mst3_arsize; initial mst3_arsize=3;

reg [2:0] slv0_awsize; initial slv0_awsize=3;
reg [2:0] slv1_awsize; initial slv1_awsize=3;
reg [2:0] slv2_awsize; initial slv2_awsize=3;
reg [2:0] slv3_awsize; initial slv3_awsize=3;
reg [2:0] slv4_awsize; initial slv4_awsize=3;
reg [2:0] slv5_awsize; initial slv5_awsize=3;
reg [2:0] slv6_awsize; initial slv6_awsize=3;
reg [2:0] slv7_awsize; initial slv7_awsize=3;
reg [2:0] slv8_awsize; initial slv8_awsize=3;
reg [2:0] slv9_awsize; initial slv9_awsize=3;
reg [2:0] slv10_awsize; initial slv10_awsize=3;
reg [2:0] slv11_awsize; initial slv11_awsize=3;
reg [2:0] slv12_awsize; initial slv12_awsize=3;
reg [2:0] slv13_awsize; initial slv13_awsize=3;
reg [2:0] slv14_awsize; initial slv14_awsize=3;
reg [2:0] slv15_awsize; initial slv15_awsize=3;

reg [2:0] slv0_arsize; initial slv0_arsize=3;
reg [2:0] slv1_arsize; initial slv1_arsize=3;
reg [2:0] slv2_arsize; initial slv2_arsize=3;
reg [2:0] slv3_arsize; initial slv3_arsize=3;
reg [2:0] slv4_arsize; initial slv4_arsize=3;
reg [2:0] slv5_arsize; initial slv5_arsize=3;
reg [2:0] slv6_arsize; initial slv6_arsize=3;
reg [2:0] slv7_arsize; initial slv7_arsize=3;
reg [2:0] slv8_arsize; initial slv8_arsize=3;
reg [2:0] slv9_arsize; initial slv9_arsize=3;
reg [2:0] slv10_arsize; initial slv10_arsize=3;
reg [2:0] slv11_arsize; initial slv11_arsize=3;
reg [2:0] slv12_arsize; initial slv12_arsize=3;
reg [2:0] slv13_arsize; initial slv13_arsize=3;
reg [2:0] slv14_arsize; initial slv14_arsize=3;
reg [2:0] slv15_arsize; initial slv15_arsize=3;

parameter IDWID = 4;
parameter DWID = 64;
parameter EXTRAS = 8;
parameter WSTRB = (DWID / 8);
reg  clk;
reg [31:0] mst0_araddr;
reg [1:0] mst0_arburst;
reg [(EXTRAS - 1):0] mst0_arextras;
reg [(IDWID - 1):0] mst0_arid;
reg [7:0] mst0_arlen;
wire  mst0_arready;
reg  mst0_arvalid;
reg [31:0] mst0_awaddr;
reg [1:0] mst0_awburst;
reg [(EXTRAS - 1):0] mst0_awextras;
reg [(IDWID - 1):0] mst0_awid;
reg [7:0] mst0_awlen;
wire  mst0_awready;
reg  mst0_awvalid;
wire [(IDWID - 1):0] mst0_bid;
reg  mst0_bready;
wire [1:0] mst0_bresp;
wire  mst0_bvalid;
wire [(DWID - 1):0] mst0_rdata;
wire [(IDWID - 1):0] mst0_rid;
wire  mst0_rlast;
reg  mst0_rready;
wire [1:0] mst0_rresp;
wire  mst0_rvalid;
reg [(DWID - 1):0] mst0_wdata;
reg  mst0_wlast;
wire  mst0_wready;
reg [(WSTRB - 1):0] mst0_wstrb;
reg  mst0_wvalid;
reg [31:0] mst1_araddr;
reg [1:0] mst1_arburst;
reg [(EXTRAS - 1):0] mst1_arextras;
reg [(IDWID - 1):0] mst1_arid;
reg [7:0] mst1_arlen;
wire  mst1_arready;
reg  mst1_arvalid;
reg [31:0] mst1_awaddr;
reg [1:0] mst1_awburst;
reg [(EXTRAS - 1):0] mst1_awextras;
reg [(IDWID - 1):0] mst1_awid;
reg [7:0] mst1_awlen;
wire  mst1_awready;
reg  mst1_awvalid;
wire [(IDWID - 1):0] mst1_bid;
reg  mst1_bready;
wire [1:0] mst1_bresp;
wire  mst1_bvalid;
wire [(DWID - 1):0] mst1_rdata;
wire [(IDWID - 1):0] mst1_rid;
wire  mst1_rlast;
reg  mst1_rready;
wire [1:0] mst1_rresp;
wire  mst1_rvalid;
reg [(DWID - 1):0] mst1_wdata;
reg  mst1_wlast;
wire  mst1_wready;
reg [(WSTRB - 1):0] mst1_wstrb;
reg  mst1_wvalid;
reg [31:0] mst2_araddr;
reg [1:0] mst2_arburst;
reg [(EXTRAS - 1):0] mst2_arextras;
reg [(IDWID - 1):0] mst2_arid;
reg [7:0] mst2_arlen;
wire  mst2_arready;
reg  mst2_arvalid;
reg [31:0] mst2_awaddr;
reg [1:0] mst2_awburst;
reg [(EXTRAS - 1):0] mst2_awextras;
reg [(IDWID - 1):0] mst2_awid;
reg [7:0] mst2_awlen;
wire  mst2_awready;
reg  mst2_awvalid;
wire [(IDWID - 1):0] mst2_bid;
reg  mst2_bready;
wire [1:0] mst2_bresp;
wire  mst2_bvalid;
wire [(DWID - 1):0] mst2_rdata;
wire [(IDWID - 1):0] mst2_rid;
wire  mst2_rlast;
reg  mst2_rready;
wire [1:0] mst2_rresp;
wire  mst2_rvalid;
reg [(DWID - 1):0] mst2_wdata;
reg  mst2_wlast;
wire  mst2_wready;
reg [(WSTRB - 1):0] mst2_wstrb;
reg  mst2_wvalid;
reg [31:0] mst3_araddr;
reg [1:0] mst3_arburst;
reg [(EXTRAS - 1):0] mst3_arextras;
reg [(IDWID - 1):0] mst3_arid;
reg [7:0] mst3_arlen;
wire  mst3_arready;
reg  mst3_arvalid;
reg [31:0] mst3_awaddr;
reg [1:0] mst3_awburst;
reg [(EXTRAS - 1):0] mst3_awextras;
reg [(IDWID - 1):0] mst3_awid;
reg [7:0] mst3_awlen;
wire  mst3_awready;
reg  mst3_awvalid;
wire [(IDWID - 1):0] mst3_bid;
reg  mst3_bready;
wire [1:0] mst3_bresp;
wire  mst3_bvalid;
wire [(DWID - 1):0] mst3_rdata;
wire [(IDWID - 1):0] mst3_rid;
wire  mst3_rlast;
reg  mst3_rready;
wire [1:0] mst3_rresp;
wire  mst3_rvalid;
reg [(DWID - 1):0] mst3_wdata;
reg  mst3_wlast;
wire  mst3_wready;
reg [(WSTRB - 1):0] mst3_wstrb;
reg  mst3_wvalid;
reg  rst_n;
wire [31:0] slv0_araddr;
wire [1:0] slv0_arburst;
wire [(EXTRAS - 1):0] slv0_arextras;
wire [(IDWID - 1):0] slv0_arid;
wire [7:0] slv0_arlen;
reg  slv0_arready;
wire  slv0_arvalid;
wire [31:0] slv0_awaddr;
wire [1:0] slv0_awburst;
wire [(EXTRAS - 1):0] slv0_awextras;
wire [(IDWID - 1):0] slv0_awid;
wire [7:0] slv0_awlen;
reg  slv0_awready;
wire  slv0_awvalid;
reg [(IDWID - 1):0] slv0_bid;
wire  slv0_bready;
reg [1:0] slv0_bresp;
reg  slv0_bvalid;
reg [(DWID - 1):0] slv0_rdata;
reg [(IDWID - 1):0] slv0_rid;
reg  slv0_rlast;
wire  slv0_rready;
reg [1:0] slv0_rresp;
reg  slv0_rvalid;
wire [(DWID - 1):0] slv0_wdata;
wire  slv0_wlast;
reg  slv0_wready;
wire [(WSTRB - 1):0] slv0_wstrb;
wire  slv0_wvalid;
wire [31:0] slv10_araddr;
wire [1:0] slv10_arburst;
wire [(EXTRAS - 1):0] slv10_arextras;
wire [(IDWID - 1):0] slv10_arid;
wire [7:0] slv10_arlen;
reg  slv10_arready;
wire  slv10_arvalid;
wire [31:0] slv10_awaddr;
wire [1:0] slv10_awburst;
wire [(EXTRAS - 1):0] slv10_awextras;
wire [(IDWID - 1):0] slv10_awid;
wire [7:0] slv10_awlen;
reg  slv10_awready;
wire  slv10_awvalid;
reg [(IDWID - 1):0] slv10_bid;
wire  slv10_bready;
reg [1:0] slv10_bresp;
reg  slv10_bvalid;
reg [(DWID - 1):0] slv10_rdata;
reg [(IDWID - 1):0] slv10_rid;
reg  slv10_rlast;
wire  slv10_rready;
reg [1:0] slv10_rresp;
reg  slv10_rvalid;
wire [(DWID - 1):0] slv10_wdata;
wire  slv10_wlast;
reg  slv10_wready;
wire [(WSTRB - 1):0] slv10_wstrb;
wire  slv10_wvalid;
wire [31:0] slv11_araddr;
wire [1:0] slv11_arburst;
wire [(EXTRAS - 1):0] slv11_arextras;
wire [(IDWID - 1):0] slv11_arid;
wire [7:0] slv11_arlen;
reg  slv11_arready;
wire  slv11_arvalid;
wire [31:0] slv11_awaddr;
wire [1:0] slv11_awburst;
wire [(EXTRAS - 1):0] slv11_awextras;
wire [(IDWID - 1):0] slv11_awid;
wire [7:0] slv11_awlen;
reg  slv11_awready;
wire  slv11_awvalid;
reg [(IDWID - 1):0] slv11_bid;
wire  slv11_bready;
reg [1:0] slv11_bresp;
reg  slv11_bvalid;
reg [(DWID - 1):0] slv11_rdata;
reg [(IDWID - 1):0] slv11_rid;
reg  slv11_rlast;
wire  slv11_rready;
reg [1:0] slv11_rresp;
reg  slv11_rvalid;
wire [(DWID - 1):0] slv11_wdata;
wire  slv11_wlast;
reg  slv11_wready;
wire [(WSTRB - 1):0] slv11_wstrb;
wire  slv11_wvalid;
wire [31:0] slv12_araddr;
wire [1:0] slv12_arburst;
wire [(EXTRAS - 1):0] slv12_arextras;
wire [(IDWID - 1):0] slv12_arid;
wire [7:0] slv12_arlen;
reg  slv12_arready;
wire  slv12_arvalid;
wire [31:0] slv12_awaddr;
wire [1:0] slv12_awburst;
wire [(EXTRAS - 1):0] slv12_awextras;
wire [(IDWID - 1):0] slv12_awid;
wire [7:0] slv12_awlen;
reg  slv12_awready;
wire  slv12_awvalid;
reg [(IDWID - 1):0] slv12_bid;
wire  slv12_bready;
reg [1:0] slv12_bresp;
reg  slv12_bvalid;
reg [(DWID - 1):0] slv12_rdata;
reg [(IDWID - 1):0] slv12_rid;
reg  slv12_rlast;
wire  slv12_rready;
reg [1:0] slv12_rresp;
reg  slv12_rvalid;
wire [(DWID - 1):0] slv12_wdata;
wire  slv12_wlast;
reg  slv12_wready;
wire [(WSTRB - 1):0] slv12_wstrb;
wire  slv12_wvalid;
wire [31:0] slv13_araddr;
wire [1:0] slv13_arburst;
wire [(EXTRAS - 1):0] slv13_arextras;
wire [(IDWID - 1):0] slv13_arid;
wire [7:0] slv13_arlen;
reg  slv13_arready;
wire  slv13_arvalid;
wire [31:0] slv13_awaddr;
wire [1:0] slv13_awburst;
wire [(EXTRAS - 1):0] slv13_awextras;
wire [(IDWID - 1):0] slv13_awid;
wire [7:0] slv13_awlen;
reg  slv13_awready;
wire  slv13_awvalid;
reg [(IDWID - 1):0] slv13_bid;
wire  slv13_bready;
reg [1:0] slv13_bresp;
reg  slv13_bvalid;
reg [(DWID - 1):0] slv13_rdata;
reg [(IDWID - 1):0] slv13_rid;
reg  slv13_rlast;
wire  slv13_rready;
reg [1:0] slv13_rresp;
reg  slv13_rvalid;
wire [(DWID - 1):0] slv13_wdata;
wire  slv13_wlast;
reg  slv13_wready;
wire [(WSTRB - 1):0] slv13_wstrb;
wire  slv13_wvalid;
wire [31:0] slv14_araddr;
wire [1:0] slv14_arburst;
wire [(EXTRAS - 1):0] slv14_arextras;
wire [(IDWID - 1):0] slv14_arid;
wire [7:0] slv14_arlen;
reg  slv14_arready;
wire  slv14_arvalid;
wire [31:0] slv14_awaddr;
wire [1:0] slv14_awburst;
wire [(EXTRAS - 1):0] slv14_awextras;
wire [(IDWID - 1):0] slv14_awid;
wire [7:0] slv14_awlen;
reg  slv14_awready;
wire  slv14_awvalid;
reg [(IDWID - 1):0] slv14_bid;
wire  slv14_bready;
reg [1:0] slv14_bresp;
reg  slv14_bvalid;
reg [(DWID - 1):0] slv14_rdata;
reg [(IDWID - 1):0] slv14_rid;
reg  slv14_rlast;
wire  slv14_rready;
reg [1:0] slv14_rresp;
reg  slv14_rvalid;
wire [(DWID - 1):0] slv14_wdata;
wire  slv14_wlast;
reg  slv14_wready;
wire [(WSTRB - 1):0] slv14_wstrb;
wire  slv14_wvalid;
wire [31:0] slv15_araddr;
wire [1:0] slv15_arburst;
wire [(EXTRAS - 1):0] slv15_arextras;
wire [(IDWID - 1):0] slv15_arid;
wire [7:0] slv15_arlen;
reg  slv15_arready;
wire  slv15_arvalid;
wire [31:0] slv15_awaddr;
wire [1:0] slv15_awburst;
wire [(EXTRAS - 1):0] slv15_awextras;
wire [(IDWID - 1):0] slv15_awid;
wire [7:0] slv15_awlen;
reg  slv15_awready;
wire  slv15_awvalid;
reg [(IDWID - 1):0] slv15_bid;
wire  slv15_bready;
reg [1:0] slv15_bresp;
reg  slv15_bvalid;
reg [(DWID - 1):0] slv15_rdata;
reg [(IDWID - 1):0] slv15_rid;
reg  slv15_rlast;
wire  slv15_rready;
reg [1:0] slv15_rresp;
reg  slv15_rvalid;
wire [(DWID - 1):0] slv15_wdata;
wire  slv15_wlast;
reg  slv15_wready;
wire [(WSTRB - 1):0] slv15_wstrb;
wire  slv15_wvalid;
wire [31:0] slv1_araddr;
wire [1:0] slv1_arburst;
wire [(EXTRAS - 1):0] slv1_arextras;
wire [(IDWID - 1):0] slv1_arid;
wire [7:0] slv1_arlen;
reg  slv1_arready;
wire  slv1_arvalid;
wire [31:0] slv1_awaddr;
wire [1:0] slv1_awburst;
wire [(EXTRAS - 1):0] slv1_awextras;
wire [(IDWID - 1):0] slv1_awid;
wire [7:0] slv1_awlen;
reg  slv1_awready;
wire  slv1_awvalid;
reg [(IDWID - 1):0] slv1_bid;
wire  slv1_bready;
reg [1:0] slv1_bresp;
reg  slv1_bvalid;
reg [(DWID - 1):0] slv1_rdata;
reg [(IDWID - 1):0] slv1_rid;
reg  slv1_rlast;
wire  slv1_rready;
reg [1:0] slv1_rresp;
reg  slv1_rvalid;
wire [(DWID - 1):0] slv1_wdata;
wire  slv1_wlast;
reg  slv1_wready;
wire [(WSTRB - 1):0] slv1_wstrb;
wire  slv1_wvalid;
wire [31:0] slv2_araddr;
wire [1:0] slv2_arburst;
wire [(EXTRAS - 1):0] slv2_arextras;
wire [(IDWID - 1):0] slv2_arid;
wire [7:0] slv2_arlen;
reg  slv2_arready;
wire  slv2_arvalid;
wire [31:0] slv2_awaddr;
wire [1:0] slv2_awburst;
wire [(EXTRAS - 1):0] slv2_awextras;
wire [(IDWID - 1):0] slv2_awid;
wire [7:0] slv2_awlen;
reg  slv2_awready;
wire  slv2_awvalid;
reg [(IDWID - 1):0] slv2_bid;
wire  slv2_bready;
reg [1:0] slv2_bresp;
reg  slv2_bvalid;
reg [(DWID - 1):0] slv2_rdata;
reg [(IDWID - 1):0] slv2_rid;
reg  slv2_rlast;
wire  slv2_rready;
reg [1:0] slv2_rresp;
reg  slv2_rvalid;
wire [(DWID - 1):0] slv2_wdata;
wire  slv2_wlast;
reg  slv2_wready;
wire [(WSTRB - 1):0] slv2_wstrb;
wire  slv2_wvalid;
wire [31:0] slv3_araddr;
wire [1:0] slv3_arburst;
wire [(EXTRAS - 1):0] slv3_arextras;
wire [(IDWID - 1):0] slv3_arid;
wire [7:0] slv3_arlen;
reg  slv3_arready;
wire  slv3_arvalid;
wire [31:0] slv3_awaddr;
wire [1:0] slv3_awburst;
wire [(EXTRAS - 1):0] slv3_awextras;
wire [(IDWID - 1):0] slv3_awid;
wire [7:0] slv3_awlen;
reg  slv3_awready;
wire  slv3_awvalid;
reg [(IDWID - 1):0] slv3_bid;
wire  slv3_bready;
reg [1:0] slv3_bresp;
reg  slv3_bvalid;
reg [(DWID - 1):0] slv3_rdata;
reg [(IDWID - 1):0] slv3_rid;
reg  slv3_rlast;
wire  slv3_rready;
reg [1:0] slv3_rresp;
reg  slv3_rvalid;
wire [(DWID - 1):0] slv3_wdata;
wire  slv3_wlast;
reg  slv3_wready;
wire [(WSTRB - 1):0] slv3_wstrb;
wire  slv3_wvalid;
wire [31:0] slv4_araddr;
wire [1:0] slv4_arburst;
wire [(EXTRAS - 1):0] slv4_arextras;
wire [(IDWID - 1):0] slv4_arid;
wire [7:0] slv4_arlen;
reg  slv4_arready;
wire  slv4_arvalid;
wire [31:0] slv4_awaddr;
wire [1:0] slv4_awburst;
wire [(EXTRAS - 1):0] slv4_awextras;
wire [(IDWID - 1):0] slv4_awid;
wire [7:0] slv4_awlen;
reg  slv4_awready;
wire  slv4_awvalid;
reg [(IDWID - 1):0] slv4_bid;
wire  slv4_bready;
reg [1:0] slv4_bresp;
reg  slv4_bvalid;
reg [(DWID - 1):0] slv4_rdata;
reg [(IDWID - 1):0] slv4_rid;
reg  slv4_rlast;
wire  slv4_rready;
reg [1:0] slv4_rresp;
reg  slv4_rvalid;
wire [(DWID - 1):0] slv4_wdata;
wire  slv4_wlast;
reg  slv4_wready;
wire [(WSTRB - 1):0] slv4_wstrb;
wire  slv4_wvalid;
wire [31:0] slv5_araddr;
wire [1:0] slv5_arburst;
wire [(EXTRAS - 1):0] slv5_arextras;
wire [(IDWID - 1):0] slv5_arid;
wire [7:0] slv5_arlen;
reg  slv5_arready;
wire  slv5_arvalid;
wire [31:0] slv5_awaddr;
wire [1:0] slv5_awburst;
wire [(EXTRAS - 1):0] slv5_awextras;
wire [(IDWID - 1):0] slv5_awid;
wire [7:0] slv5_awlen;
reg  slv5_awready;
wire  slv5_awvalid;
reg [(IDWID - 1):0] slv5_bid;
wire  slv5_bready;
reg [1:0] slv5_bresp;
reg  slv5_bvalid;
reg [(DWID - 1):0] slv5_rdata;
reg [(IDWID - 1):0] slv5_rid;
reg  slv5_rlast;
wire  slv5_rready;
reg [1:0] slv5_rresp;
reg  slv5_rvalid;
wire [(DWID - 1):0] slv5_wdata;
wire  slv5_wlast;
reg  slv5_wready;
wire [(WSTRB - 1):0] slv5_wstrb;
wire  slv5_wvalid;
wire [31:0] slv6_araddr;
wire [1:0] slv6_arburst;
wire [(EXTRAS - 1):0] slv6_arextras;
wire [(IDWID - 1):0] slv6_arid;
wire [7:0] slv6_arlen;
reg  slv6_arready;
wire  slv6_arvalid;
wire [31:0] slv6_awaddr;
wire [1:0] slv6_awburst;
wire [(EXTRAS - 1):0] slv6_awextras;
wire [(IDWID - 1):0] slv6_awid;
wire [7:0] slv6_awlen;
reg  slv6_awready;
wire  slv6_awvalid;
reg [(IDWID - 1):0] slv6_bid;
wire  slv6_bready;
reg [1:0] slv6_bresp;
reg  slv6_bvalid;
reg [(DWID - 1):0] slv6_rdata;
reg [(IDWID - 1):0] slv6_rid;
reg  slv6_rlast;
wire  slv6_rready;
reg [1:0] slv6_rresp;
reg  slv6_rvalid;
wire [(DWID - 1):0] slv6_wdata;
wire  slv6_wlast;
reg  slv6_wready;
wire [(WSTRB - 1):0] slv6_wstrb;
wire  slv6_wvalid;
wire [31:0] slv7_araddr;
wire [1:0] slv7_arburst;
wire [(EXTRAS - 1):0] slv7_arextras;
wire [(IDWID - 1):0] slv7_arid;
wire [7:0] slv7_arlen;
reg  slv7_arready;
wire  slv7_arvalid;
wire [31:0] slv7_awaddr;
wire [1:0] slv7_awburst;
wire [(EXTRAS - 1):0] slv7_awextras;
wire [(IDWID - 1):0] slv7_awid;
wire [7:0] slv7_awlen;
reg  slv7_awready;
wire  slv7_awvalid;
reg [(IDWID - 1):0] slv7_bid;
wire  slv7_bready;
reg [1:0] slv7_bresp;
reg  slv7_bvalid;
reg [(DWID - 1):0] slv7_rdata;
reg [(IDWID - 1):0] slv7_rid;
reg  slv7_rlast;
wire  slv7_rready;
reg [1:0] slv7_rresp;
reg  slv7_rvalid;
wire [(DWID - 1):0] slv7_wdata;
wire  slv7_wlast;
reg  slv7_wready;
wire [(WSTRB - 1):0] slv7_wstrb;
wire  slv7_wvalid;
wire [31:0] slv8_araddr;
wire [1:0] slv8_arburst;
wire [(EXTRAS - 1):0] slv8_arextras;
wire [(IDWID - 1):0] slv8_arid;
wire [7:0] slv8_arlen;
reg  slv8_arready;
wire  slv8_arvalid;
wire [31:0] slv8_awaddr;
wire [1:0] slv8_awburst;
wire [(EXTRAS - 1):0] slv8_awextras;
wire [(IDWID - 1):0] slv8_awid;
wire [7:0] slv8_awlen;
reg  slv8_awready;
wire  slv8_awvalid;
reg [(IDWID - 1):0] slv8_bid;
wire  slv8_bready;
reg [1:0] slv8_bresp;
reg  slv8_bvalid;
reg [(DWID - 1):0] slv8_rdata;
reg [(IDWID - 1):0] slv8_rid;
reg  slv8_rlast;
wire  slv8_rready;
reg [1:0] slv8_rresp;
reg  slv8_rvalid;
wire [(DWID - 1):0] slv8_wdata;
wire  slv8_wlast;
reg  slv8_wready;
wire [(WSTRB - 1):0] slv8_wstrb;
wire  slv8_wvalid;
wire [31:0] slv9_araddr;
wire [1:0] slv9_arburst;
wire [(EXTRAS - 1):0] slv9_arextras;
wire [(IDWID - 1):0] slv9_arid;
wire [7:0] slv9_arlen;
reg  slv9_arready;
wire  slv9_arvalid;
wire [31:0] slv9_awaddr;
wire [1:0] slv9_awburst;
wire [(EXTRAS - 1):0] slv9_awextras;
wire [(IDWID - 1):0] slv9_awid;
wire [7:0] slv9_awlen;
reg  slv9_awready;
wire  slv9_awvalid;
reg [(IDWID - 1):0] slv9_bid;
wire  slv9_bready;
reg [1:0] slv9_bresp;
reg  slv9_bvalid;
reg [(DWID - 1):0] slv9_rdata;
reg [(IDWID - 1):0] slv9_rid;
reg  slv9_rlast;
wire  slv9_rready;
reg [1:0] slv9_rresp;
reg  slv9_rvalid;
wire [(DWID - 1):0] slv9_wdata;
wire  slv9_wlast;
reg  slv9_wready;
wire [(WSTRB - 1):0] slv9_wstrb;
wire  slv9_wvalid;

always begin
    clk=0;
    #10;
    clk=1;
    #3;
    $python("negedge()");
    #7;
end
initial begin
    $dumpvars(0,tb);
    clk = 0;
    mst0_araddr = 0;
    mst0_arburst = 0;
    mst0_arextras = 0;
    mst0_arid = 0;
    mst0_arlen = 0;
    mst0_arvalid = 0;
    mst0_awaddr = 0;
    mst0_awburst = 0;
    mst0_awextras = 0;
    mst0_awid = 0;
    mst0_awlen = 0;
    mst0_awvalid = 0;
    mst0_bready = 0;
    mst0_rready = 0;
    mst0_wdata = 0;
    mst0_wlast = 0;
    mst0_wstrb = 0;
    mst0_wvalid = 0;
    mst1_araddr = 0;
    mst1_arburst = 0;
    mst1_arextras = 0;
    mst1_arid = 0;
    mst1_arlen = 0;
    mst1_arvalid = 0;
    mst1_awaddr = 0;
    mst1_awburst = 0;
    mst1_awextras = 0;
    mst1_awid = 0;
    mst1_awlen = 0;
    mst1_awvalid = 0;
    mst1_bready = 0;
    mst1_rready = 0;
    mst1_wdata = 0;
    mst1_wlast = 0;
    mst1_wstrb = 0;
    mst1_wvalid = 0;
    mst2_araddr = 0;
    mst2_arburst = 0;
    mst2_arextras = 0;
    mst2_arid = 0;
    mst2_arlen = 0;
    mst2_arvalid = 0;
    mst2_awaddr = 0;
    mst2_awburst = 0;
    mst2_awextras = 0;
    mst2_awid = 0;
    mst2_awlen = 0;
    mst2_awvalid = 0;
    mst2_bready = 0;
    mst2_rready = 0;
    mst2_wdata = 0;
    mst2_wlast = 0;
    mst2_wstrb = 0;
    mst2_wvalid = 0;
    mst3_araddr = 0;
    mst3_arburst = 0;
    mst3_arextras = 0;
    mst3_arid = 0;
    mst3_arlen = 0;
    mst3_arvalid = 0;
    mst3_awaddr = 0;
    mst3_awburst = 0;
    mst3_awextras = 0;
    mst3_awid = 0;
    mst3_awlen = 0;
    mst3_awvalid = 0;
    mst3_bready = 0;
    mst3_rready = 0;
    mst3_wdata = 0;
    mst3_wlast = 0;
    mst3_wstrb = 0;
    mst3_wvalid = 0;
    rst_n = 0;
    slv0_arready = 0;
    slv0_awready = 0;
    slv0_bid = 0;
    slv0_bresp = 0;
    slv0_bvalid = 0;
    slv0_rdata = 0;
    slv0_rid = 0;
    slv0_rlast = 0;
    slv0_rresp = 0;
    slv0_rvalid = 0;
    slv0_wready = 0;
    slv10_arready = 0;
    slv10_awready = 0;
    slv10_bid = 0;
    slv10_bresp = 0;
    slv10_bvalid = 0;
    slv10_rdata = 0;
    slv10_rid = 0;
    slv10_rlast = 0;
    slv10_rresp = 0;
    slv10_rvalid = 0;
    slv10_wready = 0;
    slv11_arready = 0;
    slv11_awready = 0;
    slv11_bid = 0;
    slv11_bresp = 0;
    slv11_bvalid = 0;
    slv11_rdata = 0;
    slv11_rid = 0;
    slv11_rlast = 0;
    slv11_rresp = 0;
    slv11_rvalid = 0;
    slv11_wready = 0;
    slv12_arready = 0;
    slv12_awready = 0;
    slv12_bid = 0;
    slv12_bresp = 0;
    slv12_bvalid = 0;
    slv12_rdata = 0;
    slv12_rid = 0;
    slv12_rlast = 0;
    slv12_rresp = 0;
    slv12_rvalid = 0;
    slv12_wready = 0;
    slv13_arready = 0;
    slv13_awready = 0;
    slv13_bid = 0;
    slv13_bresp = 0;
    slv13_bvalid = 0;
    slv13_rdata = 0;
    slv13_rid = 0;
    slv13_rlast = 0;
    slv13_rresp = 0;
    slv13_rvalid = 0;
    slv13_wready = 0;
    slv14_arready = 0;
    slv14_awready = 0;
    slv14_bid = 0;
    slv14_bresp = 0;
    slv14_bvalid = 0;
    slv14_rdata = 0;
    slv14_rid = 0;
    slv14_rlast = 0;
    slv14_rresp = 0;
    slv14_rvalid = 0;
    slv14_wready = 0;
    slv15_arready = 0;
    slv15_awready = 0;
    slv15_bid = 0;
    slv15_bresp = 0;
    slv15_bvalid = 0;
    slv15_rdata = 0;
    slv15_rid = 0;
    slv15_rlast = 0;
    slv15_rresp = 0;
    slv15_rvalid = 0;
    slv15_wready = 0;
    slv1_arready = 0;
    slv1_awready = 0;
    slv1_bid = 0;
    slv1_bresp = 0;
    slv1_bvalid = 0;
    slv1_rdata = 0;
    slv1_rid = 0;
    slv1_rlast = 0;
    slv1_rresp = 0;
    slv1_rvalid = 0;
    slv1_wready = 0;
    slv2_arready = 0;
    slv2_awready = 0;
    slv2_bid = 0;
    slv2_bresp = 0;
    slv2_bvalid = 0;
    slv2_rdata = 0;
    slv2_rid = 0;
    slv2_rlast = 0;
    slv2_rresp = 0;
    slv2_rvalid = 0;
    slv2_wready = 0;
    slv3_arready = 0;
    slv3_awready = 0;
    slv3_bid = 0;
    slv3_bresp = 0;
    slv3_bvalid = 0;
    slv3_rdata = 0;
    slv3_rid = 0;
    slv3_rlast = 0;
    slv3_rresp = 0;
    slv3_rvalid = 0;
    slv3_wready = 0;
    slv4_arready = 0;
    slv4_awready = 0;
    slv4_bid = 0;
    slv4_bresp = 0;
    slv4_bvalid = 0;
    slv4_rdata = 0;
    slv4_rid = 0;
    slv4_rlast = 0;
    slv4_rresp = 0;
    slv4_rvalid = 0;
    slv4_wready = 0;
    slv5_arready = 0;
    slv5_awready = 0;
    slv5_bid = 0;
    slv5_bresp = 0;
    slv5_bvalid = 0;
    slv5_rdata = 0;
    slv5_rid = 0;
    slv5_rlast = 0;
    slv5_rresp = 0;
    slv5_rvalid = 0;
    slv5_wready = 0;
    slv6_arready = 0;
    slv6_awready = 0;
    slv6_bid = 0;
    slv6_bresp = 0;
    slv6_bvalid = 0;
    slv6_rdata = 0;
    slv6_rid = 0;
    slv6_rlast = 0;
    slv6_rresp = 0;
    slv6_rvalid = 0;
    slv6_wready = 0;
    slv7_arready = 0;
    slv7_awready = 0;
    slv7_bid = 0;
    slv7_bresp = 0;
    slv7_bvalid = 0;
    slv7_rdata = 0;
    slv7_rid = 0;
    slv7_rlast = 0;
    slv7_rresp = 0;
    slv7_rvalid = 0;
    slv7_wready = 0;
    slv8_arready = 0;
    slv8_awready = 0;
    slv8_bid = 0;
    slv8_bresp = 0;
    slv8_bvalid = 0;
    slv8_rdata = 0;
    slv8_rid = 0;
    slv8_rlast = 0;
    slv8_rresp = 0;
    slv8_rvalid = 0;
    slv8_wready = 0;
    slv9_arready = 0;
    slv9_awready = 0;
    slv9_bid = 0;
    slv9_bresp = 0;
    slv9_bvalid = 0;
    slv9_rdata = 0;
    slv9_rid = 0;
    slv9_rlast = 0;
    slv9_rresp = 0;
    slv9_rvalid = 0;
    slv9_wready = 0;
    #100;
    rst_n=1;
end
test0 dut (
     .clk(clk)
    ,.mst0_araddr(mst0_araddr[31:0])
    ,.mst0_arburst(mst0_arburst[1:0])
    ,.mst0_arextras(mst0_arextras[(EXTRAS - 1):0])
    ,.mst0_arid(mst0_arid[(IDWID - 1):0])
    ,.mst0_arlen(mst0_arlen[7:0])
    ,.mst0_arready(mst0_arready)
    ,.mst0_arvalid(mst0_arvalid)
    ,.mst0_awaddr(mst0_awaddr[31:0])
    ,.mst0_awburst(mst0_awburst[1:0])
    ,.mst0_awextras(mst0_awextras[(EXTRAS - 1):0])
    ,.mst0_awid(mst0_awid[(IDWID - 1):0])
    ,.mst0_awlen(mst0_awlen[7:0])
    ,.mst0_awready(mst0_awready)
    ,.mst0_awvalid(mst0_awvalid)
    ,.mst0_bid(mst0_bid[(IDWID - 1):0])
    ,.mst0_bready(mst0_bready)
    ,.mst0_bresp(mst0_bresp[1:0])
    ,.mst0_bvalid(mst0_bvalid)
    ,.mst0_rdata(mst0_rdata[(DWID - 1):0])
    ,.mst0_rid(mst0_rid[(IDWID - 1):0])
    ,.mst0_rlast(mst0_rlast)
    ,.mst0_rready(mst0_rready)
    ,.mst0_rresp(mst0_rresp[1:0])
    ,.mst0_rvalid(mst0_rvalid)
    ,.mst0_wdata(mst0_wdata[(DWID - 1):0])
    ,.mst0_wlast(mst0_wlast)
    ,.mst0_wready(mst0_wready)
    ,.mst0_wstrb(mst0_wstrb[(WSTRB - 1):0])
    ,.mst0_wvalid(mst0_wvalid)
    ,.mst1_araddr(mst1_araddr[31:0])
    ,.mst1_arburst(mst1_arburst[1:0])
    ,.mst1_arextras(mst1_arextras[(EXTRAS - 1):0])
    ,.mst1_arid(mst1_arid[(IDWID - 1):0])
    ,.mst1_arlen(mst1_arlen[7:0])
    ,.mst1_arready(mst1_arready)
    ,.mst1_arvalid(mst1_arvalid)
    ,.mst1_awaddr(mst1_awaddr[31:0])
    ,.mst1_awburst(mst1_awburst[1:0])
    ,.mst1_awextras(mst1_awextras[(EXTRAS - 1):0])
    ,.mst1_awid(mst1_awid[(IDWID - 1):0])
    ,.mst1_awlen(mst1_awlen[7:0])
    ,.mst1_awready(mst1_awready)
    ,.mst1_awvalid(mst1_awvalid)
    ,.mst1_bid(mst1_bid[(IDWID - 1):0])
    ,.mst1_bready(mst1_bready)
    ,.mst1_bresp(mst1_bresp[1:0])
    ,.mst1_bvalid(mst1_bvalid)
    ,.mst1_rdata(mst1_rdata[(DWID - 1):0])
    ,.mst1_rid(mst1_rid[(IDWID - 1):0])
    ,.mst1_rlast(mst1_rlast)
    ,.mst1_rready(mst1_rready)
    ,.mst1_rresp(mst1_rresp[1:0])
    ,.mst1_rvalid(mst1_rvalid)
    ,.mst1_wdata(mst1_wdata[(DWID - 1):0])
    ,.mst1_wlast(mst1_wlast)
    ,.mst1_wready(mst1_wready)
    ,.mst1_wstrb(mst1_wstrb[(WSTRB - 1):0])
    ,.mst1_wvalid(mst1_wvalid)
    ,.mst2_araddr(mst2_araddr[31:0])
    ,.mst2_arburst(mst2_arburst[1:0])
    ,.mst2_arextras(mst2_arextras[(EXTRAS - 1):0])
    ,.mst2_arid(mst2_arid[(IDWID - 1):0])
    ,.mst2_arlen(mst2_arlen[7:0])
    ,.mst2_arready(mst2_arready)
    ,.mst2_arvalid(mst2_arvalid)
    ,.mst2_awaddr(mst2_awaddr[31:0])
    ,.mst2_awburst(mst2_awburst[1:0])
    ,.mst2_awextras(mst2_awextras[(EXTRAS - 1):0])
    ,.mst2_awid(mst2_awid[(IDWID - 1):0])
    ,.mst2_awlen(mst2_awlen[7:0])
    ,.mst2_awready(mst2_awready)
    ,.mst2_awvalid(mst2_awvalid)
    ,.mst2_bid(mst2_bid[(IDWID - 1):0])
    ,.mst2_bready(mst2_bready)
    ,.mst2_bresp(mst2_bresp[1:0])
    ,.mst2_bvalid(mst2_bvalid)
    ,.mst2_rdata(mst2_rdata[(DWID - 1):0])
    ,.mst2_rid(mst2_rid[(IDWID - 1):0])
    ,.mst2_rlast(mst2_rlast)
    ,.mst2_rready(mst2_rready)
    ,.mst2_rresp(mst2_rresp[1:0])
    ,.mst2_rvalid(mst2_rvalid)
    ,.mst2_wdata(mst2_wdata[(DWID - 1):0])
    ,.mst2_wlast(mst2_wlast)
    ,.mst2_wready(mst2_wready)
    ,.mst2_wstrb(mst2_wstrb[(WSTRB - 1):0])
    ,.mst2_wvalid(mst2_wvalid)
    ,.mst3_araddr(mst3_araddr[31:0])
    ,.mst3_arburst(mst3_arburst[1:0])
    ,.mst3_arextras(mst3_arextras[(EXTRAS - 1):0])
    ,.mst3_arid(mst3_arid[(IDWID - 1):0])
    ,.mst3_arlen(mst3_arlen[7:0])
    ,.mst3_arready(mst3_arready)
    ,.mst3_arvalid(mst3_arvalid)
    ,.mst3_awaddr(mst3_awaddr[31:0])
    ,.mst3_awburst(mst3_awburst[1:0])
    ,.mst3_awextras(mst3_awextras[(EXTRAS - 1):0])
    ,.mst3_awid(mst3_awid[(IDWID - 1):0])
    ,.mst3_awlen(mst3_awlen[7:0])
    ,.mst3_awready(mst3_awready)
    ,.mst3_awvalid(mst3_awvalid)
    ,.mst3_bid(mst3_bid[(IDWID - 1):0])
    ,.mst3_bready(mst3_bready)
    ,.mst3_bresp(mst3_bresp[1:0])
    ,.mst3_bvalid(mst3_bvalid)
    ,.mst3_rdata(mst3_rdata[(DWID - 1):0])
    ,.mst3_rid(mst3_rid[(IDWID - 1):0])
    ,.mst3_rlast(mst3_rlast)
    ,.mst3_rready(mst3_rready)
    ,.mst3_rresp(mst3_rresp[1:0])
    ,.mst3_rvalid(mst3_rvalid)
    ,.mst3_wdata(mst3_wdata[(DWID - 1):0])
    ,.mst3_wlast(mst3_wlast)
    ,.mst3_wready(mst3_wready)
    ,.mst3_wstrb(mst3_wstrb[(WSTRB - 1):0])
    ,.mst3_wvalid(mst3_wvalid)
    ,.rst_n(rst_n)
    ,.slv0_araddr(slv0_araddr[31:0])
    ,.slv0_arburst(slv0_arburst[1:0])
    ,.slv0_arextras(slv0_arextras[(EXTRAS - 1):0])
    ,.slv0_arid(slv0_arid[(IDWID - 1):0])
    ,.slv0_arlen(slv0_arlen[7:0])
    ,.slv0_arready(slv0_arready)
    ,.slv0_arvalid(slv0_arvalid)
    ,.slv0_awaddr(slv0_awaddr[31:0])
    ,.slv0_awburst(slv0_awburst[1:0])
    ,.slv0_awextras(slv0_awextras[(EXTRAS - 1):0])
    ,.slv0_awid(slv0_awid[(IDWID - 1):0])
    ,.slv0_awlen(slv0_awlen[7:0])
    ,.slv0_awready(slv0_awready)
    ,.slv0_awvalid(slv0_awvalid)
    ,.slv0_bid(slv0_bid[(IDWID - 1):0])
    ,.slv0_bready(slv0_bready)
    ,.slv0_bresp(slv0_bresp[1:0])
    ,.slv0_bvalid(slv0_bvalid)
    ,.slv0_rdata(slv0_rdata[(DWID - 1):0])
    ,.slv0_rid(slv0_rid[(IDWID - 1):0])
    ,.slv0_rlast(slv0_rlast)
    ,.slv0_rready(slv0_rready)
    ,.slv0_rresp(slv0_rresp[1:0])
    ,.slv0_rvalid(slv0_rvalid)
    ,.slv0_wdata(slv0_wdata[(DWID - 1):0])
    ,.slv0_wlast(slv0_wlast)
    ,.slv0_wready(slv0_wready)
    ,.slv0_wstrb(slv0_wstrb[(WSTRB - 1):0])
    ,.slv0_wvalid(slv0_wvalid)
    ,.slv10_araddr(slv10_araddr[31:0])
    ,.slv10_arburst(slv10_arburst[1:0])
    ,.slv10_arextras(slv10_arextras[(EXTRAS - 1):0])
    ,.slv10_arid(slv10_arid[(IDWID - 1):0])
    ,.slv10_arlen(slv10_arlen[7:0])
    ,.slv10_arready(slv10_arready)
    ,.slv10_arvalid(slv10_arvalid)
    ,.slv10_awaddr(slv10_awaddr[31:0])
    ,.slv10_awburst(slv10_awburst[1:0])
    ,.slv10_awextras(slv10_awextras[(EXTRAS - 1):0])
    ,.slv10_awid(slv10_awid[(IDWID - 1):0])
    ,.slv10_awlen(slv10_awlen[7:0])
    ,.slv10_awready(slv10_awready)
    ,.slv10_awvalid(slv10_awvalid)
    ,.slv10_bid(slv10_bid[(IDWID - 1):0])
    ,.slv10_bready(slv10_bready)
    ,.slv10_bresp(slv10_bresp[1:0])
    ,.slv10_bvalid(slv10_bvalid)
    ,.slv10_rdata(slv10_rdata[(DWID - 1):0])
    ,.slv10_rid(slv10_rid[(IDWID - 1):0])
    ,.slv10_rlast(slv10_rlast)
    ,.slv10_rready(slv10_rready)
    ,.slv10_rresp(slv10_rresp[1:0])
    ,.slv10_rvalid(slv10_rvalid)
    ,.slv10_wdata(slv10_wdata[(DWID - 1):0])
    ,.slv10_wlast(slv10_wlast)
    ,.slv10_wready(slv10_wready)
    ,.slv10_wstrb(slv10_wstrb[(WSTRB - 1):0])
    ,.slv10_wvalid(slv10_wvalid)
    ,.slv11_araddr(slv11_araddr[31:0])
    ,.slv11_arburst(slv11_arburst[1:0])
    ,.slv11_arextras(slv11_arextras[(EXTRAS - 1):0])
    ,.slv11_arid(slv11_arid[(IDWID - 1):0])
    ,.slv11_arlen(slv11_arlen[7:0])
    ,.slv11_arready(slv11_arready)
    ,.slv11_arvalid(slv11_arvalid)
    ,.slv11_awaddr(slv11_awaddr[31:0])
    ,.slv11_awburst(slv11_awburst[1:0])
    ,.slv11_awextras(slv11_awextras[(EXTRAS - 1):0])
    ,.slv11_awid(slv11_awid[(IDWID - 1):0])
    ,.slv11_awlen(slv11_awlen[7:0])
    ,.slv11_awready(slv11_awready)
    ,.slv11_awvalid(slv11_awvalid)
    ,.slv11_bid(slv11_bid[(IDWID - 1):0])
    ,.slv11_bready(slv11_bready)
    ,.slv11_bresp(slv11_bresp[1:0])
    ,.slv11_bvalid(slv11_bvalid)
    ,.slv11_rdata(slv11_rdata[(DWID - 1):0])
    ,.slv11_rid(slv11_rid[(IDWID - 1):0])
    ,.slv11_rlast(slv11_rlast)
    ,.slv11_rready(slv11_rready)
    ,.slv11_rresp(slv11_rresp[1:0])
    ,.slv11_rvalid(slv11_rvalid)
    ,.slv11_wdata(slv11_wdata[(DWID - 1):0])
    ,.slv11_wlast(slv11_wlast)
    ,.slv11_wready(slv11_wready)
    ,.slv11_wstrb(slv11_wstrb[(WSTRB - 1):0])
    ,.slv11_wvalid(slv11_wvalid)
    ,.slv12_araddr(slv12_araddr[31:0])
    ,.slv12_arburst(slv12_arburst[1:0])
    ,.slv12_arextras(slv12_arextras[(EXTRAS - 1):0])
    ,.slv12_arid(slv12_arid[(IDWID - 1):0])
    ,.slv12_arlen(slv12_arlen[7:0])
    ,.slv12_arready(slv12_arready)
    ,.slv12_arvalid(slv12_arvalid)
    ,.slv12_awaddr(slv12_awaddr[31:0])
    ,.slv12_awburst(slv12_awburst[1:0])
    ,.slv12_awextras(slv12_awextras[(EXTRAS - 1):0])
    ,.slv12_awid(slv12_awid[(IDWID - 1):0])
    ,.slv12_awlen(slv12_awlen[7:0])
    ,.slv12_awready(slv12_awready)
    ,.slv12_awvalid(slv12_awvalid)
    ,.slv12_bid(slv12_bid[(IDWID - 1):0])
    ,.slv12_bready(slv12_bready)
    ,.slv12_bresp(slv12_bresp[1:0])
    ,.slv12_bvalid(slv12_bvalid)
    ,.slv12_rdata(slv12_rdata[(DWID - 1):0])
    ,.slv12_rid(slv12_rid[(IDWID - 1):0])
    ,.slv12_rlast(slv12_rlast)
    ,.slv12_rready(slv12_rready)
    ,.slv12_rresp(slv12_rresp[1:0])
    ,.slv12_rvalid(slv12_rvalid)
    ,.slv12_wdata(slv12_wdata[(DWID - 1):0])
    ,.slv12_wlast(slv12_wlast)
    ,.slv12_wready(slv12_wready)
    ,.slv12_wstrb(slv12_wstrb[(WSTRB - 1):0])
    ,.slv12_wvalid(slv12_wvalid)
    ,.slv13_araddr(slv13_araddr[31:0])
    ,.slv13_arburst(slv13_arburst[1:0])
    ,.slv13_arextras(slv13_arextras[(EXTRAS - 1):0])
    ,.slv13_arid(slv13_arid[(IDWID - 1):0])
    ,.slv13_arlen(slv13_arlen[7:0])
    ,.slv13_arready(slv13_arready)
    ,.slv13_arvalid(slv13_arvalid)
    ,.slv13_awaddr(slv13_awaddr[31:0])
    ,.slv13_awburst(slv13_awburst[1:0])
    ,.slv13_awextras(slv13_awextras[(EXTRAS - 1):0])
    ,.slv13_awid(slv13_awid[(IDWID - 1):0])
    ,.slv13_awlen(slv13_awlen[7:0])
    ,.slv13_awready(slv13_awready)
    ,.slv13_awvalid(slv13_awvalid)
    ,.slv13_bid(slv13_bid[(IDWID - 1):0])
    ,.slv13_bready(slv13_bready)
    ,.slv13_bresp(slv13_bresp[1:0])
    ,.slv13_bvalid(slv13_bvalid)
    ,.slv13_rdata(slv13_rdata[(DWID - 1):0])
    ,.slv13_rid(slv13_rid[(IDWID - 1):0])
    ,.slv13_rlast(slv13_rlast)
    ,.slv13_rready(slv13_rready)
    ,.slv13_rresp(slv13_rresp[1:0])
    ,.slv13_rvalid(slv13_rvalid)
    ,.slv13_wdata(slv13_wdata[(DWID - 1):0])
    ,.slv13_wlast(slv13_wlast)
    ,.slv13_wready(slv13_wready)
    ,.slv13_wstrb(slv13_wstrb[(WSTRB - 1):0])
    ,.slv13_wvalid(slv13_wvalid)
    ,.slv14_araddr(slv14_araddr[31:0])
    ,.slv14_arburst(slv14_arburst[1:0])
    ,.slv14_arextras(slv14_arextras[(EXTRAS - 1):0])
    ,.slv14_arid(slv14_arid[(IDWID - 1):0])
    ,.slv14_arlen(slv14_arlen[7:0])
    ,.slv14_arready(slv14_arready)
    ,.slv14_arvalid(slv14_arvalid)
    ,.slv14_awaddr(slv14_awaddr[31:0])
    ,.slv14_awburst(slv14_awburst[1:0])
    ,.slv14_awextras(slv14_awextras[(EXTRAS - 1):0])
    ,.slv14_awid(slv14_awid[(IDWID - 1):0])
    ,.slv14_awlen(slv14_awlen[7:0])
    ,.slv14_awready(slv14_awready)
    ,.slv14_awvalid(slv14_awvalid)
    ,.slv14_bid(slv14_bid[(IDWID - 1):0])
    ,.slv14_bready(slv14_bready)
    ,.slv14_bresp(slv14_bresp[1:0])
    ,.slv14_bvalid(slv14_bvalid)
    ,.slv14_rdata(slv14_rdata[(DWID - 1):0])
    ,.slv14_rid(slv14_rid[(IDWID - 1):0])
    ,.slv14_rlast(slv14_rlast)
    ,.slv14_rready(slv14_rready)
    ,.slv14_rresp(slv14_rresp[1:0])
    ,.slv14_rvalid(slv14_rvalid)
    ,.slv14_wdata(slv14_wdata[(DWID - 1):0])
    ,.slv14_wlast(slv14_wlast)
    ,.slv14_wready(slv14_wready)
    ,.slv14_wstrb(slv14_wstrb[(WSTRB - 1):0])
    ,.slv14_wvalid(slv14_wvalid)
    ,.slv15_araddr(slv15_araddr[31:0])
    ,.slv15_arburst(slv15_arburst[1:0])
    ,.slv15_arextras(slv15_arextras[(EXTRAS - 1):0])
    ,.slv15_arid(slv15_arid[(IDWID - 1):0])
    ,.slv15_arlen(slv15_arlen[7:0])
    ,.slv15_arready(slv15_arready)
    ,.slv15_arvalid(slv15_arvalid)
    ,.slv15_awaddr(slv15_awaddr[31:0])
    ,.slv15_awburst(slv15_awburst[1:0])
    ,.slv15_awextras(slv15_awextras[(EXTRAS - 1):0])
    ,.slv15_awid(slv15_awid[(IDWID - 1):0])
    ,.slv15_awlen(slv15_awlen[7:0])
    ,.slv15_awready(slv15_awready)
    ,.slv15_awvalid(slv15_awvalid)
    ,.slv15_bid(slv15_bid[(IDWID - 1):0])
    ,.slv15_bready(slv15_bready)
    ,.slv15_bresp(slv15_bresp[1:0])
    ,.slv15_bvalid(slv15_bvalid)
    ,.slv15_rdata(slv15_rdata[(DWID - 1):0])
    ,.slv15_rid(slv15_rid[(IDWID - 1):0])
    ,.slv15_rlast(slv15_rlast)
    ,.slv15_rready(slv15_rready)
    ,.slv15_rresp(slv15_rresp[1:0])
    ,.slv15_rvalid(slv15_rvalid)
    ,.slv15_wdata(slv15_wdata[(DWID - 1):0])
    ,.slv15_wlast(slv15_wlast)
    ,.slv15_wready(slv15_wready)
    ,.slv15_wstrb(slv15_wstrb[(WSTRB - 1):0])
    ,.slv15_wvalid(slv15_wvalid)
    ,.slv1_araddr(slv1_araddr[31:0])
    ,.slv1_arburst(slv1_arburst[1:0])
    ,.slv1_arextras(slv1_arextras[(EXTRAS - 1):0])
    ,.slv1_arid(slv1_arid[(IDWID - 1):0])
    ,.slv1_arlen(slv1_arlen[7:0])
    ,.slv1_arready(slv1_arready)
    ,.slv1_arvalid(slv1_arvalid)
    ,.slv1_awaddr(slv1_awaddr[31:0])
    ,.slv1_awburst(slv1_awburst[1:0])
    ,.slv1_awextras(slv1_awextras[(EXTRAS - 1):0])
    ,.slv1_awid(slv1_awid[(IDWID - 1):0])
    ,.slv1_awlen(slv1_awlen[7:0])
    ,.slv1_awready(slv1_awready)
    ,.slv1_awvalid(slv1_awvalid)
    ,.slv1_bid(slv1_bid[(IDWID - 1):0])
    ,.slv1_bready(slv1_bready)
    ,.slv1_bresp(slv1_bresp[1:0])
    ,.slv1_bvalid(slv1_bvalid)
    ,.slv1_rdata(slv1_rdata[(DWID - 1):0])
    ,.slv1_rid(slv1_rid[(IDWID - 1):0])
    ,.slv1_rlast(slv1_rlast)
    ,.slv1_rready(slv1_rready)
    ,.slv1_rresp(slv1_rresp[1:0])
    ,.slv1_rvalid(slv1_rvalid)
    ,.slv1_wdata(slv1_wdata[(DWID - 1):0])
    ,.slv1_wlast(slv1_wlast)
    ,.slv1_wready(slv1_wready)
    ,.slv1_wstrb(slv1_wstrb[(WSTRB - 1):0])
    ,.slv1_wvalid(slv1_wvalid)
    ,.slv2_araddr(slv2_araddr[31:0])
    ,.slv2_arburst(slv2_arburst[1:0])
    ,.slv2_arextras(slv2_arextras[(EXTRAS - 1):0])
    ,.slv2_arid(slv2_arid[(IDWID - 1):0])
    ,.slv2_arlen(slv2_arlen[7:0])
    ,.slv2_arready(slv2_arready)
    ,.slv2_arvalid(slv2_arvalid)
    ,.slv2_awaddr(slv2_awaddr[31:0])
    ,.slv2_awburst(slv2_awburst[1:0])
    ,.slv2_awextras(slv2_awextras[(EXTRAS - 1):0])
    ,.slv2_awid(slv2_awid[(IDWID - 1):0])
    ,.slv2_awlen(slv2_awlen[7:0])
    ,.slv2_awready(slv2_awready)
    ,.slv2_awvalid(slv2_awvalid)
    ,.slv2_bid(slv2_bid[(IDWID - 1):0])
    ,.slv2_bready(slv2_bready)
    ,.slv2_bresp(slv2_bresp[1:0])
    ,.slv2_bvalid(slv2_bvalid)
    ,.slv2_rdata(slv2_rdata[(DWID - 1):0])
    ,.slv2_rid(slv2_rid[(IDWID - 1):0])
    ,.slv2_rlast(slv2_rlast)
    ,.slv2_rready(slv2_rready)
    ,.slv2_rresp(slv2_rresp[1:0])
    ,.slv2_rvalid(slv2_rvalid)
    ,.slv2_wdata(slv2_wdata[(DWID - 1):0])
    ,.slv2_wlast(slv2_wlast)
    ,.slv2_wready(slv2_wready)
    ,.slv2_wstrb(slv2_wstrb[(WSTRB - 1):0])
    ,.slv2_wvalid(slv2_wvalid)
    ,.slv3_araddr(slv3_araddr[31:0])
    ,.slv3_arburst(slv3_arburst[1:0])
    ,.slv3_arextras(slv3_arextras[(EXTRAS - 1):0])
    ,.slv3_arid(slv3_arid[(IDWID - 1):0])
    ,.slv3_arlen(slv3_arlen[7:0])
    ,.slv3_arready(slv3_arready)
    ,.slv3_arvalid(slv3_arvalid)
    ,.slv3_awaddr(slv3_awaddr[31:0])
    ,.slv3_awburst(slv3_awburst[1:0])
    ,.slv3_awextras(slv3_awextras[(EXTRAS - 1):0])
    ,.slv3_awid(slv3_awid[(IDWID - 1):0])
    ,.slv3_awlen(slv3_awlen[7:0])
    ,.slv3_awready(slv3_awready)
    ,.slv3_awvalid(slv3_awvalid)
    ,.slv3_bid(slv3_bid[(IDWID - 1):0])
    ,.slv3_bready(slv3_bready)
    ,.slv3_bresp(slv3_bresp[1:0])
    ,.slv3_bvalid(slv3_bvalid)
    ,.slv3_rdata(slv3_rdata[(DWID - 1):0])
    ,.slv3_rid(slv3_rid[(IDWID - 1):0])
    ,.slv3_rlast(slv3_rlast)
    ,.slv3_rready(slv3_rready)
    ,.slv3_rresp(slv3_rresp[1:0])
    ,.slv3_rvalid(slv3_rvalid)
    ,.slv3_wdata(slv3_wdata[(DWID - 1):0])
    ,.slv3_wlast(slv3_wlast)
    ,.slv3_wready(slv3_wready)
    ,.slv3_wstrb(slv3_wstrb[(WSTRB - 1):0])
    ,.slv3_wvalid(slv3_wvalid)
    ,.slv4_araddr(slv4_araddr[31:0])
    ,.slv4_arburst(slv4_arburst[1:0])
    ,.slv4_arextras(slv4_arextras[(EXTRAS - 1):0])
    ,.slv4_arid(slv4_arid[(IDWID - 1):0])
    ,.slv4_arlen(slv4_arlen[7:0])
    ,.slv4_arready(slv4_arready)
    ,.slv4_arvalid(slv4_arvalid)
    ,.slv4_awaddr(slv4_awaddr[31:0])
    ,.slv4_awburst(slv4_awburst[1:0])
    ,.slv4_awextras(slv4_awextras[(EXTRAS - 1):0])
    ,.slv4_awid(slv4_awid[(IDWID - 1):0])
    ,.slv4_awlen(slv4_awlen[7:0])
    ,.slv4_awready(slv4_awready)
    ,.slv4_awvalid(slv4_awvalid)
    ,.slv4_bid(slv4_bid[(IDWID - 1):0])
    ,.slv4_bready(slv4_bready)
    ,.slv4_bresp(slv4_bresp[1:0])
    ,.slv4_bvalid(slv4_bvalid)
    ,.slv4_rdata(slv4_rdata[(DWID - 1):0])
    ,.slv4_rid(slv4_rid[(IDWID - 1):0])
    ,.slv4_rlast(slv4_rlast)
    ,.slv4_rready(slv4_rready)
    ,.slv4_rresp(slv4_rresp[1:0])
    ,.slv4_rvalid(slv4_rvalid)
    ,.slv4_wdata(slv4_wdata[(DWID - 1):0])
    ,.slv4_wlast(slv4_wlast)
    ,.slv4_wready(slv4_wready)
    ,.slv4_wstrb(slv4_wstrb[(WSTRB - 1):0])
    ,.slv4_wvalid(slv4_wvalid)
    ,.slv5_araddr(slv5_araddr[31:0])
    ,.slv5_arburst(slv5_arburst[1:0])
    ,.slv5_arextras(slv5_arextras[(EXTRAS - 1):0])
    ,.slv5_arid(slv5_arid[(IDWID - 1):0])
    ,.slv5_arlen(slv5_arlen[7:0])
    ,.slv5_arready(slv5_arready)
    ,.slv5_arvalid(slv5_arvalid)
    ,.slv5_awaddr(slv5_awaddr[31:0])
    ,.slv5_awburst(slv5_awburst[1:0])
    ,.slv5_awextras(slv5_awextras[(EXTRAS - 1):0])
    ,.slv5_awid(slv5_awid[(IDWID - 1):0])
    ,.slv5_awlen(slv5_awlen[7:0])
    ,.slv5_awready(slv5_awready)
    ,.slv5_awvalid(slv5_awvalid)
    ,.slv5_bid(slv5_bid[(IDWID - 1):0])
    ,.slv5_bready(slv5_bready)
    ,.slv5_bresp(slv5_bresp[1:0])
    ,.slv5_bvalid(slv5_bvalid)
    ,.slv5_rdata(slv5_rdata[(DWID - 1):0])
    ,.slv5_rid(slv5_rid[(IDWID - 1):0])
    ,.slv5_rlast(slv5_rlast)
    ,.slv5_rready(slv5_rready)
    ,.slv5_rresp(slv5_rresp[1:0])
    ,.slv5_rvalid(slv5_rvalid)
    ,.slv5_wdata(slv5_wdata[(DWID - 1):0])
    ,.slv5_wlast(slv5_wlast)
    ,.slv5_wready(slv5_wready)
    ,.slv5_wstrb(slv5_wstrb[(WSTRB - 1):0])
    ,.slv5_wvalid(slv5_wvalid)
    ,.slv6_araddr(slv6_araddr[31:0])
    ,.slv6_arburst(slv6_arburst[1:0])
    ,.slv6_arextras(slv6_arextras[(EXTRAS - 1):0])
    ,.slv6_arid(slv6_arid[(IDWID - 1):0])
    ,.slv6_arlen(slv6_arlen[7:0])
    ,.slv6_arready(slv6_arready)
    ,.slv6_arvalid(slv6_arvalid)
    ,.slv6_awaddr(slv6_awaddr[31:0])
    ,.slv6_awburst(slv6_awburst[1:0])
    ,.slv6_awextras(slv6_awextras[(EXTRAS - 1):0])
    ,.slv6_awid(slv6_awid[(IDWID - 1):0])
    ,.slv6_awlen(slv6_awlen[7:0])
    ,.slv6_awready(slv6_awready)
    ,.slv6_awvalid(slv6_awvalid)
    ,.slv6_bid(slv6_bid[(IDWID - 1):0])
    ,.slv6_bready(slv6_bready)
    ,.slv6_bresp(slv6_bresp[1:0])
    ,.slv6_bvalid(slv6_bvalid)
    ,.slv6_rdata(slv6_rdata[(DWID - 1):0])
    ,.slv6_rid(slv6_rid[(IDWID - 1):0])
    ,.slv6_rlast(slv6_rlast)
    ,.slv6_rready(slv6_rready)
    ,.slv6_rresp(slv6_rresp[1:0])
    ,.slv6_rvalid(slv6_rvalid)
    ,.slv6_wdata(slv6_wdata[(DWID - 1):0])
    ,.slv6_wlast(slv6_wlast)
    ,.slv6_wready(slv6_wready)
    ,.slv6_wstrb(slv6_wstrb[(WSTRB - 1):0])
    ,.slv6_wvalid(slv6_wvalid)
    ,.slv7_araddr(slv7_araddr[31:0])
    ,.slv7_arburst(slv7_arburst[1:0])
    ,.slv7_arextras(slv7_arextras[(EXTRAS - 1):0])
    ,.slv7_arid(slv7_arid[(IDWID - 1):0])
    ,.slv7_arlen(slv7_arlen[7:0])
    ,.slv7_arready(slv7_arready)
    ,.slv7_arvalid(slv7_arvalid)
    ,.slv7_awaddr(slv7_awaddr[31:0])
    ,.slv7_awburst(slv7_awburst[1:0])
    ,.slv7_awextras(slv7_awextras[(EXTRAS - 1):0])
    ,.slv7_awid(slv7_awid[(IDWID - 1):0])
    ,.slv7_awlen(slv7_awlen[7:0])
    ,.slv7_awready(slv7_awready)
    ,.slv7_awvalid(slv7_awvalid)
    ,.slv7_bid(slv7_bid[(IDWID - 1):0])
    ,.slv7_bready(slv7_bready)
    ,.slv7_bresp(slv7_bresp[1:0])
    ,.slv7_bvalid(slv7_bvalid)
    ,.slv7_rdata(slv7_rdata[(DWID - 1):0])
    ,.slv7_rid(slv7_rid[(IDWID - 1):0])
    ,.slv7_rlast(slv7_rlast)
    ,.slv7_rready(slv7_rready)
    ,.slv7_rresp(slv7_rresp[1:0])
    ,.slv7_rvalid(slv7_rvalid)
    ,.slv7_wdata(slv7_wdata[(DWID - 1):0])
    ,.slv7_wlast(slv7_wlast)
    ,.slv7_wready(slv7_wready)
    ,.slv7_wstrb(slv7_wstrb[(WSTRB - 1):0])
    ,.slv7_wvalid(slv7_wvalid)
    ,.slv8_araddr(slv8_araddr[31:0])
    ,.slv8_arburst(slv8_arburst[1:0])
    ,.slv8_arextras(slv8_arextras[(EXTRAS - 1):0])
    ,.slv8_arid(slv8_arid[(IDWID - 1):0])
    ,.slv8_arlen(slv8_arlen[7:0])
    ,.slv8_arready(slv8_arready)
    ,.slv8_arvalid(slv8_arvalid)
    ,.slv8_awaddr(slv8_awaddr[31:0])
    ,.slv8_awburst(slv8_awburst[1:0])
    ,.slv8_awextras(slv8_awextras[(EXTRAS - 1):0])
    ,.slv8_awid(slv8_awid[(IDWID - 1):0])
    ,.slv8_awlen(slv8_awlen[7:0])
    ,.slv8_awready(slv8_awready)
    ,.slv8_awvalid(slv8_awvalid)
    ,.slv8_bid(slv8_bid[(IDWID - 1):0])
    ,.slv8_bready(slv8_bready)
    ,.slv8_bresp(slv8_bresp[1:0])
    ,.slv8_bvalid(slv8_bvalid)
    ,.slv8_rdata(slv8_rdata[(DWID - 1):0])
    ,.slv8_rid(slv8_rid[(IDWID - 1):0])
    ,.slv8_rlast(slv8_rlast)
    ,.slv8_rready(slv8_rready)
    ,.slv8_rresp(slv8_rresp[1:0])
    ,.slv8_rvalid(slv8_rvalid)
    ,.slv8_wdata(slv8_wdata[(DWID - 1):0])
    ,.slv8_wlast(slv8_wlast)
    ,.slv8_wready(slv8_wready)
    ,.slv8_wstrb(slv8_wstrb[(WSTRB - 1):0])
    ,.slv8_wvalid(slv8_wvalid)
    ,.slv9_araddr(slv9_araddr[31:0])
    ,.slv9_arburst(slv9_arburst[1:0])
    ,.slv9_arextras(slv9_arextras[(EXTRAS - 1):0])
    ,.slv9_arid(slv9_arid[(IDWID - 1):0])
    ,.slv9_arlen(slv9_arlen[7:0])
    ,.slv9_arready(slv9_arready)
    ,.slv9_arvalid(slv9_arvalid)
    ,.slv9_awaddr(slv9_awaddr[31:0])
    ,.slv9_awburst(slv9_awburst[1:0])
    ,.slv9_awextras(slv9_awextras[(EXTRAS - 1):0])
    ,.slv9_awid(slv9_awid[(IDWID - 1):0])
    ,.slv9_awlen(slv9_awlen[7:0])
    ,.slv9_awready(slv9_awready)
    ,.slv9_awvalid(slv9_awvalid)
    ,.slv9_bid(slv9_bid[(IDWID - 1):0])
    ,.slv9_bready(slv9_bready)
    ,.slv9_bresp(slv9_bresp[1:0])
    ,.slv9_bvalid(slv9_bvalid)
    ,.slv9_rdata(slv9_rdata[(DWID - 1):0])
    ,.slv9_rid(slv9_rid[(IDWID - 1):0])
    ,.slv9_rlast(slv9_rlast)
    ,.slv9_rready(slv9_rready)
    ,.slv9_rresp(slv9_rresp[1:0])
    ,.slv9_rvalid(slv9_rvalid)
    ,.slv9_wdata(slv9_wdata[(DWID - 1):0])
    ,.slv9_wlast(slv9_wlast)
    ,.slv9_wready(slv9_wready)
    ,.slv9_wstrb(slv9_wstrb[(WSTRB - 1):0])
    ,.slv9_wvalid(slv9_wvalid)
);

reg [1023:0] testname;
initial begin
   if ($value$plusargs("LOG=%s",testname)) begin 
        $python("pymonname()",testname);
    end 


    if ($value$plusargs("SEQ=%s",testname)) begin 
         $display(" Running SEQ= %s.",testname); 
    end else begin
        testname = 0;
        $display(" default test");
    end 
    #10;
    if (testname!=0) $python("sequence()",testname);
end 
endmodule

