module atan_table_till_10(input [9:0] addr,output [24:0] result,output [24:0] lastone);
assign result = 
    (addr==0) ? 18574873 :  //   in=2.000000 val=1.107149
    (addr==1) ? 18601005 :  //   in=2.007812 val=1.108706
    (addr==2) ? 18626976 :  //   in=2.015625 val=1.110254
    (addr==3) ? 18652785 :  //   in=2.023438 val=1.111793
    (addr==4) ? 18678434 :  //   in=2.031250 val=1.113321
    (addr==5) ? 18703926 :  //   in=2.039062 val=1.114841
    (addr==6) ? 18729260 :  //   in=2.046875 val=1.116351
    (addr==7) ? 18754438 :  //   in=2.054688 val=1.117852
    (addr==8) ? 18779463 :  //   in=2.062500 val=1.119343
    (addr==9) ? 18804334 :  //   in=2.070312 val=1.120826
    (addr==10) ? 18829053 :  //   in=2.078125 val=1.122299
    (addr==11) ? 18853623 :  //   in=2.085938 val=1.123764
    (addr==12) ? 18878042 :  //   in=2.093750 val=1.125219
    (addr==13) ? 18902314 :  //   in=2.101562 val=1.126666
    (addr==14) ? 18926440 :  //   in=2.109375 val=1.128104
    (addr==15) ? 18950419 :  //   in=2.117188 val=1.129533
    (addr==16) ? 18974255 :  //   in=2.125000 val=1.130954
    (addr==17) ? 18997947 :  //   in=2.132812 val=1.132366
    (addr==18) ? 19021498 :  //   in=2.140625 val=1.133770
    (addr==19) ? 19044908 :  //   in=2.148438 val=1.135165
    (addr==20) ? 19068178 :  //   in=2.156250 val=1.136552
    (addr==21) ? 19091310 :  //   in=2.164062 val=1.137931
    (addr==22) ? 19114305 :  //   in=2.171875 val=1.139301
    (addr==23) ? 19137163 :  //   in=2.179688 val=1.140664
    (addr==24) ? 19159887 :  //   in=2.187500 val=1.142018
    (addr==25) ? 19182477 :  //   in=2.195312 val=1.143365
    (addr==26) ? 19204934 :  //   in=2.203125 val=1.144703
    (addr==27) ? 19227260 :  //   in=2.210938 val=1.146034
    (addr==28) ? 19249454 :  //   in=2.218750 val=1.147357
    (addr==29) ? 19271520 :  //   in=2.226562 val=1.148672
    (addr==30) ? 19293456 :  //   in=2.234375 val=1.149980
    (addr==31) ? 19315266 :  //   in=2.242188 val=1.151280
    (addr==32) ? 19336949 :  //   in=2.250000 val=1.152572
    (addr==33) ? 19358506 :  //   in=2.257812 val=1.153857
    (addr==34) ? 19379940 :  //   in=2.265625 val=1.155134
    (addr==35) ? 19401250 :  //   in=2.273438 val=1.156405
    (addr==36) ? 19422437 :  //   in=2.281250 val=1.157667
    (addr==37) ? 19443503 :  //   in=2.289062 val=1.158923
    (addr==38) ? 19464449 :  //   in=2.296875 val=1.160172
    (addr==39) ? 19485275 :  //   in=2.304688 val=1.161413
    (addr==40) ? 19505983 :  //   in=2.312500 val=1.162647
    (addr==41) ? 19526573 :  //   in=2.320312 val=1.163874
    (addr==42) ? 19547047 :  //   in=2.328125 val=1.165095
    (addr==43) ? 19567405 :  //   in=2.335938 val=1.166308
    (addr==44) ? 19587648 :  //   in=2.343750 val=1.167515
    (addr==45) ? 19607778 :  //   in=2.351562 val=1.168715
    (addr==46) ? 19627794 :  //   in=2.359375 val=1.169908
    (addr==47) ? 19647698 :  //   in=2.367188 val=1.171094
    (addr==48) ? 19667492 :  //   in=2.375000 val=1.172274
    (addr==49) ? 19687175 :  //   in=2.382812 val=1.173447
    (addr==50) ? 19706748 :  //   in=2.390625 val=1.174614
    (addr==51) ? 19726213 :  //   in=2.398438 val=1.175774
    (addr==52) ? 19745570 :  //   in=2.406250 val=1.176928
    (addr==53) ? 19764820 :  //   in=2.414062 val=1.178075
    (addr==54) ? 19783964 :  //   in=2.421875 val=1.179216
    (addr==55) ? 19803003 :  //   in=2.429688 val=1.180351
    (addr==56) ? 19821938 :  //   in=2.437500 val=1.181480
    (addr==57) ? 19840769 :  //   in=2.445312 val=1.182602
    (addr==58) ? 19859497 :  //   in=2.453125 val=1.183718
    (addr==59) ? 19878123 :  //   in=2.460938 val=1.184829
    (addr==60) ? 19896648 :  //   in=2.468750 val=1.185933
    (addr==61) ? 19915073 :  //   in=2.476562 val=1.187031
    (addr==62) ? 19933397 :  //   in=2.484375 val=1.188123
    (addr==63) ? 19951623 :  //   in=2.492188 val=1.189209
    (addr==64) ? 19969751 :  //   in=2.500000 val=1.190290
    (addr==65) ? 19987781 :  //   in=2.507812 val=1.191365
    (addr==66) ? 20005715 :  //   in=2.515625 val=1.192434
    (addr==67) ? 20023553 :  //   in=2.523438 val=1.193497
    (addr==68) ? 20041295 :  //   in=2.531250 val=1.194554
    (addr==69) ? 20058943 :  //   in=2.539062 val=1.195606
    (addr==70) ? 20076498 :  //   in=2.546875 val=1.196653
    (addr==71) ? 20093959 :  //   in=2.554688 val=1.197693
    (addr==72) ? 20111328 :  //   in=2.562500 val=1.198729
    (addr==73) ? 20128605 :  //   in=2.570312 val=1.199758
    (addr==74) ? 20145791 :  //   in=2.578125 val=1.200783
    (addr==75) ? 20162887 :  //   in=2.585938 val=1.201802
    (addr==76) ? 20179893 :  //   in=2.593750 val=1.202815
    (addr==77) ? 20196810 :  //   in=2.601562 val=1.203824
    (addr==78) ? 20213639 :  //   in=2.609375 val=1.204827
    (addr==79) ? 20230381 :  //   in=2.617188 val=1.205825
    (addr==80) ? 20247035 :  //   in=2.625000 val=1.206817
    (addr==81) ? 20263603 :  //   in=2.632812 val=1.207805
    (addr==82) ? 20280086 :  //   in=2.640625 val=1.208787
    (addr==83) ? 20296483 :  //   in=2.648438 val=1.209765
    (addr==84) ? 20312796 :  //   in=2.656250 val=1.210737
    (addr==85) ? 20329025 :  //   in=2.664062 val=1.211704
    (addr==86) ? 20345170 :  //   in=2.671875 val=1.212667
    (addr==87) ? 20361234 :  //   in=2.679688 val=1.213624
    (addr==88) ? 20377215 :  //   in=2.687500 val=1.214577
    (addr==89) ? 20393114 :  //   in=2.695312 val=1.215524
    (addr==90) ? 20408933 :  //   in=2.703125 val=1.216467
    (addr==91) ? 20424672 :  //   in=2.710938 val=1.217405
    (addr==92) ? 20440331 :  //   in=2.718750 val=1.218339
    (addr==93) ? 20455911 :  //   in=2.726562 val=1.219267
    (addr==94) ? 20471413 :  //   in=2.734375 val=1.220191
    (addr==95) ? 20486836 :  //   in=2.742188 val=1.221111
    (addr==96) ? 20502182 :  //   in=2.750000 val=1.222025
    (addr==97) ? 20517452 :  //   in=2.757812 val=1.222935
    (addr==98) ? 20532645 :  //   in=2.765625 val=1.223841
    (addr==99) ? 20547762 :  //   in=2.773438 val=1.224742
    (addr==100) ? 20562804 :  //   in=2.781250 val=1.225639
    (addr==101) ? 20577772 :  //   in=2.789062 val=1.226531
    (addr==102) ? 20592665 :  //   in=2.796875 val=1.227419
    (addr==103) ? 20607485 :  //   in=2.804688 val=1.228302
    (addr==104) ? 20622232 :  //   in=2.812500 val=1.229181
    (addr==105) ? 20636906 :  //   in=2.820312 val=1.230055
    (addr==106) ? 20651508 :  //   in=2.828125 val=1.230926
    (addr==107) ? 20666039 :  //   in=2.835938 val=1.231792
    (addr==108) ? 20680499 :  //   in=2.843750 val=1.232654
    (addr==109) ? 20694888 :  //   in=2.851562 val=1.233511
    (addr==110) ? 20709207 :  //   in=2.859375 val=1.234365
    (addr==111) ? 20723456 :  //   in=2.867188 val=1.235214
    (addr==112) ? 20737637 :  //   in=2.875000 val=1.236059
    (addr==113) ? 20751748 :  //   in=2.882812 val=1.236901
    (addr==114) ? 20765792 :  //   in=2.890625 val=1.237738
    (addr==115) ? 20779768 :  //   in=2.898438 val=1.238571
    (addr==116) ? 20793677 :  //   in=2.906250 val=1.239400
    (addr==117) ? 20807519 :  //   in=2.914062 val=1.240225
    (addr==118) ? 20821295 :  //   in=2.921875 val=1.241046
    (addr==119) ? 20835006 :  //   in=2.929688 val=1.241863
    (addr==120) ? 20848650 :  //   in=2.937500 val=1.242676
    (addr==121) ? 20862230 :  //   in=2.945312 val=1.243486
    (addr==122) ? 20875746 :  //   in=2.953125 val=1.244291
    (addr==123) ? 20889197 :  //   in=2.960938 val=1.245093
    (addr==124) ? 20902585 :  //   in=2.968750 val=1.245891
    (addr==125) ? 20915910 :  //   in=2.976562 val=1.246685
    (addr==126) ? 20929172 :  //   in=2.984375 val=1.247476
    (addr==127) ? 20942372 :  //   in=2.992188 val=1.248263
    (addr==128) ? 20955510 :  //   in=3.000000 val=1.249046
    (addr==129) ? 20968587 :  //   in=3.007812 val=1.249825
    (addr==130) ? 20981602 :  //   in=3.015625 val=1.250601
    (addr==131) ? 20994557 :  //   in=3.023438 val=1.251373
    (addr==132) ? 21007452 :  //   in=3.031250 val=1.252142
    (addr==133) ? 21020287 :  //   in=3.039062 val=1.252907
    (addr==134) ? 21033062 :  //   in=3.046875 val=1.253668
    (addr==135) ? 21045779 :  //   in=3.054688 val=1.254426
    (addr==136) ? 21058437 :  //   in=3.062500 val=1.255181
    (addr==137) ? 21071036 :  //   in=3.070312 val=1.255932
    (addr==138) ? 21083578 :  //   in=3.078125 val=1.256679
    (addr==139) ? 21096062 :  //   in=3.085938 val=1.257423
    (addr==140) ? 21108490 :  //   in=3.093750 val=1.258164
    (addr==141) ? 21120860 :  //   in=3.101562 val=1.258901
    (addr==142) ? 21133175 :  //   in=3.109375 val=1.259635
    (addr==143) ? 21145433 :  //   in=3.117188 val=1.260366
    (addr==144) ? 21157636 :  //   in=3.125000 val=1.261093
    (addr==145) ? 21169783 :  //   in=3.132812 val=1.261817
    (addr==146) ? 21181876 :  //   in=3.140625 val=1.262538
    (addr==147) ? 21193914 :  //   in=3.148438 val=1.263256
    (addr==148) ? 21205898 :  //   in=3.156250 val=1.263970
    (addr==149) ? 21217828 :  //   in=3.164062 val=1.264681
    (addr==150) ? 21229705 :  //   in=3.171875 val=1.265389
    (addr==151) ? 21241528 :  //   in=3.179688 val=1.266094
    (addr==152) ? 21253299 :  //   in=3.187500 val=1.266795
    (addr==153) ? 21265018 :  //   in=3.195312 val=1.267494
    (addr==154) ? 21276684 :  //   in=3.203125 val=1.268189
    (addr==155) ? 21288299 :  //   in=3.210938 val=1.268882
    (addr==156) ? 21299862 :  //   in=3.218750 val=1.269571
    (addr==157) ? 21311374 :  //   in=3.226562 val=1.270257
    (addr==158) ? 21322836 :  //   in=3.234375 val=1.270940
    (addr==159) ? 21334247 :  //   in=3.242188 val=1.271620
    (addr==160) ? 21345608 :  //   in=3.250000 val=1.272297
    (addr==161) ? 21356919 :  //   in=3.257812 val=1.272972
    (addr==162) ? 21368180 :  //   in=3.265625 val=1.273643
    (addr==163) ? 21379393 :  //   in=3.273438 val=1.274311
    (addr==164) ? 21390557 :  //   in=3.281250 val=1.274977
    (addr==165) ? 21401672 :  //   in=3.289062 val=1.275639
    (addr==166) ? 21412739 :  //   in=3.296875 val=1.276299
    (addr==167) ? 21423758 :  //   in=3.304688 val=1.276955
    (addr==168) ? 21434729 :  //   in=3.312500 val=1.277609
    (addr==169) ? 21445653 :  //   in=3.320312 val=1.278261
    (addr==170) ? 21456530 :  //   in=3.328125 val=1.278909
    (addr==171) ? 21467360 :  //   in=3.335938 val=1.279554
    (addr==172) ? 21478144 :  //   in=3.343750 val=1.280197
    (addr==173) ? 21488881 :  //   in=3.351562 val=1.280837
    (addr==174) ? 21499573 :  //   in=3.359375 val=1.281474
    (addr==175) ? 21510219 :  //   in=3.367188 val=1.282109
    (addr==176) ? 21520820 :  //   in=3.375000 val=1.282741
    (addr==177) ? 21531376 :  //   in=3.382812 val=1.283370
    (addr==178) ? 21541887 :  //   in=3.390625 val=1.283997
    (addr==179) ? 21552354 :  //   in=3.398438 val=1.284620
    (addr==180) ? 21562776 :  //   in=3.406250 val=1.285242
    (addr==181) ? 21573155 :  //   in=3.414062 val=1.285860
    (addr==182) ? 21583490 :  //   in=3.421875 val=1.286476
    (addr==183) ? 21593781 :  //   in=3.429688 val=1.287090
    (addr==184) ? 21604030 :  //   in=3.437500 val=1.287701
    (addr==185) ? 21614235 :  //   in=3.445312 val=1.288309
    (addr==186) ? 21624398 :  //   in=3.453125 val=1.288915
    (addr==187) ? 21634519 :  //   in=3.460938 val=1.289518
    (addr==188) ? 21644597 :  //   in=3.468750 val=1.290119
    (addr==189) ? 21654634 :  //   in=3.476562 val=1.290717
    (addr==190) ? 21664629 :  //   in=3.484375 val=1.291313
    (addr==191) ? 21674583 :  //   in=3.492188 val=1.291906
    (addr==192) ? 21684495 :  //   in=3.500000 val=1.292497
    (addr==193) ? 21694367 :  //   in=3.507812 val=1.293085
    (addr==194) ? 21704198 :  //   in=3.515625 val=1.293671
    (addr==195) ? 21713989 :  //   in=3.523438 val=1.294255
    (addr==196) ? 21723740 :  //   in=3.531250 val=1.294836
    (addr==197) ? 21733451 :  //   in=3.539062 val=1.295415
    (addr==198) ? 21743122 :  //   in=3.546875 val=1.295991
    (addr==199) ? 21752754 :  //   in=3.554688 val=1.296565
    (addr==200) ? 21762347 :  //   in=3.562500 val=1.297137
    (addr==201) ? 21771901 :  //   in=3.570312 val=1.297706
    (addr==202) ? 21781416 :  //   in=3.578125 val=1.298274
    (addr==203) ? 21790893 :  //   in=3.585938 val=1.298838
    (addr==204) ? 21800332 :  //   in=3.593750 val=1.299401
    (addr==205) ? 21809732 :  //   in=3.601562 val=1.299961
    (addr==206) ? 21819095 :  //   in=3.609375 val=1.300519
    (addr==207) ? 21828420 :  //   in=3.617188 val=1.301075
    (addr==208) ? 21837708 :  //   in=3.625000 val=1.301629
    (addr==209) ? 21846958 :  //   in=3.632812 val=1.302180
    (addr==210) ? 21856172 :  //   in=3.640625 val=1.302729
    (addr==211) ? 21865349 :  //   in=3.648438 val=1.303276
    (addr==212) ? 21874490 :  //   in=3.656250 val=1.303821
    (addr==213) ? 21883594 :  //   in=3.664062 val=1.304364
    (addr==214) ? 21892662 :  //   in=3.671875 val=1.304904
    (addr==215) ? 21901694 :  //   in=3.679688 val=1.305443
    (addr==216) ? 21910691 :  //   in=3.687500 val=1.305979
    (addr==217) ? 21919653 :  //   in=3.695312 val=1.306513
    (addr==218) ? 21928579 :  //   in=3.703125 val=1.307045
    (addr==219) ? 21937470 :  //   in=3.710938 val=1.307575
    (addr==220) ? 21946326 :  //   in=3.718750 val=1.308103
    (addr==221) ? 21955147 :  //   in=3.726562 val=1.308629
    (addr==222) ? 21963934 :  //   in=3.734375 val=1.309153
    (addr==223) ? 21972687 :  //   in=3.742188 val=1.309674
    (addr==224) ? 21981406 :  //   in=3.750000 val=1.310194
    (addr==225) ? 21990091 :  //   in=3.757812 val=1.310712
    (addr==226) ? 21998742 :  //   in=3.765625 val=1.311227
    (addr==227) ? 22007360 :  //   in=3.773438 val=1.311741
    (addr==228) ? 22015945 :  //   in=3.781250 val=1.312253
    (addr==229) ? 22024496 :  //   in=3.789062 val=1.312762
    (addr==230) ? 22033015 :  //   in=3.796875 val=1.313270
    (addr==231) ? 22041501 :  //   in=3.804688 val=1.313776
    (addr==232) ? 22049954 :  //   in=3.812500 val=1.314280
    (addr==233) ? 22058375 :  //   in=3.820312 val=1.314782
    (addr==234) ? 22066764 :  //   in=3.828125 val=1.315282
    (addr==235) ? 22075121 :  //   in=3.835938 val=1.315780
    (addr==236) ? 22083446 :  //   in=3.843750 val=1.316276
    (addr==237) ? 22091739 :  //   in=3.851562 val=1.316770
    (addr==238) ? 22100001 :  //   in=3.859375 val=1.317263
    (addr==239) ? 22108232 :  //   in=3.867188 val=1.317753
    (addr==240) ? 22116431 :  //   in=3.875000 val=1.318242
    (addr==241) ? 22124600 :  //   in=3.882812 val=1.318729
    (addr==242) ? 22132737 :  //   in=3.890625 val=1.319214
    (addr==243) ? 22140845 :  //   in=3.898438 val=1.319697
    (addr==244) ? 22148921 :  //   in=3.906250 val=1.320179
    (addr==245) ? 22156968 :  //   in=3.914062 val=1.320658
    (addr==246) ? 22164984 :  //   in=3.921875 val=1.321136
    (addr==247) ? 22172971 :  //   in=3.929688 val=1.321612
    (addr==248) ? 22180928 :  //   in=3.937500 val=1.322086
    (addr==249) ? 22188855 :  //   in=3.945312 val=1.322559
    (addr==250) ? 22196752 :  //   in=3.953125 val=1.323030
    (addr==251) ? 22204621 :  //   in=3.960938 val=1.323499
    (addr==252) ? 22212460 :  //   in=3.968750 val=1.323966
    (addr==253) ? 22220270 :  //   in=3.976562 val=1.324431
    (addr==254) ? 22228052 :  //   in=3.984375 val=1.324895
    (addr==255) ? 22235805 :  //   in=3.992188 val=1.325357
    (addr==256) ? 22243529 :  //   in=4.000000 val=1.325818
    (addr==257) ? 22251225 :  //   in=4.007812 val=1.326276
    (addr==258) ? 22258893 :  //   in=4.015625 val=1.326733
    (addr==259) ? 22266532 :  //   in=4.023438 val=1.327189
    (addr==260) ? 22274144 :  //   in=4.031250 val=1.327642
    (addr==261) ? 22281728 :  //   in=4.039062 val=1.328095
    (addr==262) ? 22289285 :  //   in=4.046875 val=1.328545
    (addr==263) ? 22296814 :  //   in=4.054688 val=1.328994
    (addr==264) ? 22304316 :  //   in=4.062500 val=1.329441
    (addr==265) ? 22311790 :  //   in=4.070312 val=1.329886
    (addr==266) ? 22319238 :  //   in=4.078125 val=1.330330
    (addr==267) ? 22326658 :  //   in=4.085938 val=1.330773
    (addr==268) ? 22334052 :  //   in=4.093750 val=1.331213
    (addr==269) ? 22341420 :  //   in=4.101562 val=1.331652
    (addr==270) ? 22348761 :  //   in=4.109375 val=1.332090
    (addr==271) ? 22356076 :  //   in=4.117188 val=1.332526
    (addr==272) ? 22363364 :  //   in=4.125000 val=1.332960
    (addr==273) ? 22370627 :  //   in=4.132812 val=1.333393
    (addr==274) ? 22377863 :  //   in=4.140625 val=1.333825
    (addr==275) ? 22385074 :  //   in=4.148438 val=1.334254
    (addr==276) ? 22392259 :  //   in=4.156250 val=1.334683
    (addr==277) ? 22399419 :  //   in=4.164062 val=1.335109
    (addr==278) ? 22406553 :  //   in=4.171875 val=1.335535
    (addr==279) ? 22413662 :  //   in=4.179688 val=1.335958
    (addr==280) ? 22420746 :  //   in=4.187500 val=1.336381
    (addr==281) ? 22427805 :  //   in=4.195312 val=1.336801
    (addr==282) ? 22434840 :  //   in=4.203125 val=1.337221
    (addr==283) ? 22441849 :  //   in=4.210938 val=1.337638
    (addr==284) ? 22448834 :  //   in=4.218750 val=1.338055
    (addr==285) ? 22455795 :  //   in=4.226562 val=1.338470
    (addr==286) ? 22462731 :  //   in=4.234375 val=1.338883
    (addr==287) ? 22469643 :  //   in=4.242188 val=1.339295
    (addr==288) ? 22476531 :  //   in=4.250000 val=1.339706
    (addr==289) ? 22483395 :  //   in=4.257812 val=1.340115
    (addr==290) ? 22490235 :  //   in=4.265625 val=1.340522
    (addr==291) ? 22497051 :  //   in=4.273438 val=1.340929
    (addr==292) ? 22503844 :  //   in=4.281250 val=1.341334
    (addr==293) ? 22510613 :  //   in=4.289062 val=1.341737
    (addr==294) ? 22517359 :  //   in=4.296875 val=1.342139
    (addr==295) ? 22524082 :  //   in=4.304688 val=1.342540
    (addr==296) ? 22530782 :  //   in=4.312500 val=1.342939
    (addr==297) ? 22537459 :  //   in=4.320312 val=1.343337
    (addr==298) ? 22544112 :  //   in=4.328125 val=1.343734
    (addr==299) ? 22550743 :  //   in=4.335938 val=1.344129
    (addr==300) ? 22557352 :  //   in=4.343750 val=1.344523
    (addr==301) ? 22563938 :  //   in=4.351562 val=1.344916
    (addr==302) ? 22570501 :  //   in=4.359375 val=1.345307
    (addr==303) ? 22577042 :  //   in=4.367188 val=1.345697
    (addr==304) ? 22583561 :  //   in=4.375000 val=1.346085
    (addr==305) ? 22590058 :  //   in=4.382812 val=1.346472
    (addr==306) ? 22596533 :  //   in=4.390625 val=1.346858
    (addr==307) ? 22602986 :  //   in=4.398438 val=1.347243
    (addr==308) ? 22609417 :  //   in=4.406250 val=1.347626
    (addr==309) ? 22615826 :  //   in=4.414062 val=1.348008
    (addr==310) ? 22622214 :  //   in=4.421875 val=1.348389
    (addr==311) ? 22628581 :  //   in=4.429688 val=1.348769
    (addr==312) ? 22634926 :  //   in=4.437500 val=1.349147
    (addr==313) ? 22641250 :  //   in=4.445312 val=1.349524
    (addr==314) ? 22647553 :  //   in=4.453125 val=1.349899
    (addr==315) ? 22653835 :  //   in=4.460938 val=1.350274
    (addr==316) ? 22660096 :  //   in=4.468750 val=1.350647
    (addr==317) ? 22666336 :  //   in=4.476562 val=1.351019
    (addr==318) ? 22672555 :  //   in=4.484375 val=1.351390
    (addr==319) ? 22678754 :  //   in=4.492188 val=1.351759
    (addr==320) ? 22684933 :  //   in=4.500000 val=1.352127
    (addr==321) ? 22691091 :  //   in=4.507812 val=1.352494
    (addr==322) ? 22697228 :  //   in=4.515625 val=1.352860
    (addr==323) ? 22703346 :  //   in=4.523438 val=1.353225
    (addr==324) ? 22709443 :  //   in=4.531250 val=1.353588
    (addr==325) ? 22715520 :  //   in=4.539062 val=1.353951
    (addr==326) ? 22721577 :  //   in=4.546875 val=1.354312
    (addr==327) ? 22727615 :  //   in=4.554688 val=1.354671
    (addr==328) ? 22733633 :  //   in=4.562500 val=1.355030
    (addr==329) ? 22739631 :  //   in=4.570312 val=1.355388
    (addr==330) ? 22745609 :  //   in=4.578125 val=1.355744
    (addr==331) ? 22751569 :  //   in=4.585938 val=1.356099
    (addr==332) ? 22757508 :  //   in=4.593750 val=1.356453
    (addr==333) ? 22763429 :  //   in=4.601562 val=1.356806
    (addr==334) ? 22769330 :  //   in=4.609375 val=1.357158
    (addr==335) ? 22775213 :  //   in=4.617188 val=1.357508
    (addr==336) ? 22781076 :  //   in=4.625000 val=1.357858
    (addr==337) ? 22786921 :  //   in=4.632812 val=1.358206
    (addr==338) ? 22792746 :  //   in=4.640625 val=1.358554
    (addr==339) ? 22798553 :  //   in=4.648438 val=1.358900
    (addr==340) ? 22804341 :  //   in=4.656250 val=1.359245
    (addr==341) ? 22810111 :  //   in=4.664062 val=1.359589
    (addr==342) ? 22815862 :  //   in=4.671875 val=1.359931
    (addr==343) ? 22821595 :  //   in=4.679688 val=1.360273
    (addr==344) ? 22827310 :  //   in=4.687500 val=1.360614
    (addr==345) ? 22833007 :  //   in=4.695312 val=1.360953
    (addr==346) ? 22838685 :  //   in=4.703125 val=1.361292
    (addr==347) ? 22844345 :  //   in=4.710938 val=1.361629
    (addr==348) ? 22849988 :  //   in=4.718750 val=1.361965
    (addr==349) ? 22855612 :  //   in=4.726562 val=1.362301
    (addr==350) ? 22861219 :  //   in=4.734375 val=1.362635
    (addr==351) ? 22866808 :  //   in=4.742188 val=1.362968
    (addr==352) ? 22872380 :  //   in=4.750000 val=1.363300
    (addr==353) ? 22877934 :  //   in=4.757812 val=1.363631
    (addr==354) ? 22883470 :  //   in=4.765625 val=1.363961
    (addr==355) ? 22888989 :  //   in=4.773438 val=1.364290
    (addr==356) ? 22894491 :  //   in=4.781250 val=1.364618
    (addr==357) ? 22899976 :  //   in=4.789062 val=1.364945
    (addr==358) ? 22905444 :  //   in=4.796875 val=1.365271
    (addr==359) ? 22910894 :  //   in=4.804688 val=1.365596
    (addr==360) ? 22916328 :  //   in=4.812500 val=1.365920
    (addr==361) ? 22921745 :  //   in=4.820312 val=1.366242
    (addr==362) ? 22927144 :  //   in=4.828125 val=1.366564
    (addr==363) ? 22932528 :  //   in=4.835938 val=1.366885
    (addr==364) ? 22937894 :  //   in=4.843750 val=1.367205
    (addr==365) ? 22943244 :  //   in=4.851562 val=1.367524
    (addr==366) ? 22948577 :  //   in=4.859375 val=1.367842
    (addr==367) ? 22953894 :  //   in=4.867188 val=1.368159
    (addr==368) ? 22959195 :  //   in=4.875000 val=1.368475
    (addr==369) ? 22964479 :  //   in=4.882812 val=1.368790
    (addr==370) ? 22969748 :  //   in=4.890625 val=1.369104
    (addr==371) ? 22975000 :  //   in=4.898438 val=1.369417
    (addr==372) ? 22980236 :  //   in=4.906250 val=1.369729
    (addr==373) ? 22985456 :  //   in=4.914062 val=1.370040
    (addr==374) ? 22990660 :  //   in=4.921875 val=1.370350
    (addr==375) ? 22995848 :  //   in=4.929688 val=1.370659
    (addr==376) ? 23001020 :  //   in=4.937500 val=1.370968
    (addr==377) ? 23006177 :  //   in=4.945312 val=1.371275
    (addr==378) ? 23011318 :  //   in=4.953125 val=1.371581
    (addr==379) ? 23016444 :  //   in=4.960938 val=1.371887
    (addr==380) ? 23021554 :  //   in=4.968750 val=1.372192
    (addr==381) ? 23026649 :  //   in=4.976562 val=1.372495
    (addr==382) ? 23031728 :  //   in=4.984375 val=1.372798
    (addr==383) ? 23036792 :  //   in=4.992188 val=1.373100
    (addr==384) ? 23041841 :  //   in=5.000000 val=1.373401
    (addr==385) ? 23046874 :  //   in=5.007812 val=1.373701
    (addr==386) ? 23051893 :  //   in=5.015625 val=1.374000
    (addr==387) ? 23056897 :  //   in=5.023438 val=1.374298
    (addr==388) ? 23061885 :  //   in=5.031250 val=1.374596
    (addr==389) ? 23066859 :  //   in=5.039062 val=1.374892
    (addr==390) ? 23071818 :  //   in=5.046875 val=1.375188
    (addr==391) ? 23076762 :  //   in=5.054688 val=1.375482
    (addr==392) ? 23081692 :  //   in=5.062500 val=1.375776
    (addr==393) ? 23086606 :  //   in=5.070312 val=1.376069
    (addr==394) ? 23091507 :  //   in=5.078125 val=1.376361
    (addr==395) ? 23096393 :  //   in=5.085938 val=1.376652
    (addr==396) ? 23101264 :  //   in=5.093750 val=1.376943
    (addr==397) ? 23106121 :  //   in=5.101562 val=1.377232
    (addr==398) ? 23110964 :  //   in=5.109375 val=1.377521
    (addr==399) ? 23115792 :  //   in=5.117188 val=1.377809
    (addr==400) ? 23120607 :  //   in=5.125000 val=1.378096
    (addr==401) ? 23125407 :  //   in=5.132812 val=1.378382
    (addr==402) ? 23130193 :  //   in=5.140625 val=1.378667
    (addr==403) ? 23134965 :  //   in=5.148438 val=1.378951
    (addr==404) ? 23139723 :  //   in=5.156250 val=1.379235
    (addr==405) ? 23144467 :  //   in=5.164062 val=1.379518
    (addr==406) ? 23149198 :  //   in=5.171875 val=1.379800
    (addr==407) ? 23153915 :  //   in=5.179688 val=1.380081
    (addr==408) ? 23158618 :  //   in=5.187500 val=1.380361
    (addr==409) ? 23163307 :  //   in=5.195312 val=1.380641
    (addr==410) ? 23167983 :  //   in=5.203125 val=1.380919
    (addr==411) ? 23172645 :  //   in=5.210938 val=1.381197
    (addr==412) ? 23177294 :  //   in=5.218750 val=1.381474
    (addr==413) ? 23181929 :  //   in=5.226562 val=1.381751
    (addr==414) ? 23186552 :  //   in=5.234375 val=1.382026
    (addr==415) ? 23191160 :  //   in=5.242188 val=1.382301
    (addr==416) ? 23195756 :  //   in=5.250000 val=1.382575
    (addr==417) ? 23200338 :  //   in=5.257812 val=1.382848
    (addr==418) ? 23204908 :  //   in=5.265625 val=1.383120
    (addr==419) ? 23209464 :  //   in=5.273438 val=1.383392
    (addr==420) ? 23214007 :  //   in=5.281250 val=1.383663
    (addr==421) ? 23218537 :  //   in=5.289062 val=1.383933
    (addr==422) ? 23223054 :  //   in=5.296875 val=1.384202
    (addr==423) ? 23227559 :  //   in=5.304688 val=1.384470
    (addr==424) ? 23232051 :  //   in=5.312500 val=1.384738
    (addr==425) ? 23236529 :  //   in=5.320312 val=1.385005
    (addr==426) ? 23240996 :  //   in=5.328125 val=1.385271
    (addr==427) ? 23245449 :  //   in=5.335938 val=1.385537
    (addr==428) ? 23249890 :  //   in=5.343750 val=1.385801
    (addr==429) ? 23254319 :  //   in=5.351562 val=1.386065
    (addr==430) ? 23258735 :  //   in=5.359375 val=1.386329
    (addr==431) ? 23263138 :  //   in=5.367188 val=1.386591
    (addr==432) ? 23267530 :  //   in=5.375000 val=1.386853
    (addr==433) ? 23271909 :  //   in=5.382812 val=1.387114
    (addr==434) ? 23276275 :  //   in=5.390625 val=1.387374
    (addr==435) ? 23280630 :  //   in=5.398438 val=1.387634
    (addr==436) ? 23284972 :  //   in=5.406250 val=1.387893
    (addr==437) ? 23289302 :  //   in=5.414062 val=1.388151
    (addr==438) ? 23293620 :  //   in=5.421875 val=1.388408
    (addr==439) ? 23297926 :  //   in=5.429688 val=1.388665
    (addr==440) ? 23302220 :  //   in=5.437500 val=1.388921
    (addr==441) ? 23306502 :  //   in=5.445312 val=1.389176
    (addr==442) ? 23310773 :  //   in=5.453125 val=1.389430
    (addr==443) ? 23315031 :  //   in=5.460938 val=1.389684
    (addr==444) ? 23319278 :  //   in=5.468750 val=1.389937
    (addr==445) ? 23323513 :  //   in=5.476562 val=1.390190
    (addr==446) ? 23327736 :  //   in=5.484375 val=1.390441
    (addr==447) ? 23331948 :  //   in=5.492188 val=1.390692
    (addr==448) ? 23336148 :  //   in=5.500000 val=1.390943
    (addr==449) ? 23340336 :  //   in=5.507812 val=1.391192
    (addr==450) ? 23344513 :  //   in=5.515625 val=1.391441
    (addr==451) ? 23348679 :  //   in=5.523438 val=1.391690
    (addr==452) ? 23352833 :  //   in=5.531250 val=1.391937
    (addr==453) ? 23356976 :  //   in=5.539062 val=1.392184
    (addr==454) ? 23361108 :  //   in=5.546875 val=1.392431
    (addr==455) ? 23365228 :  //   in=5.554688 val=1.392676
    (addr==456) ? 23369337 :  //   in=5.562500 val=1.392921
    (addr==457) ? 23373435 :  //   in=5.570312 val=1.393165
    (addr==458) ? 23377522 :  //   in=5.578125 val=1.393409
    (addr==459) ? 23381598 :  //   in=5.585938 val=1.393652
    (addr==460) ? 23385662 :  //   in=5.593750 val=1.393894
    (addr==461) ? 23389716 :  //   in=5.601562 val=1.394136
    (addr==462) ? 23393759 :  //   in=5.609375 val=1.394377
    (addr==463) ? 23397791 :  //   in=5.617188 val=1.394617
    (addr==464) ? 23401812 :  //   in=5.625000 val=1.394857
    (addr==465) ? 23405822 :  //   in=5.632812 val=1.395096
    (addr==466) ? 23409821 :  //   in=5.640625 val=1.395334
    (addr==467) ? 23413810 :  //   in=5.648438 val=1.395572
    (addr==468) ? 23417788 :  //   in=5.656250 val=1.395809
    (addr==469) ? 23421755 :  //   in=5.664062 val=1.396045
    (addr==470) ? 23425712 :  //   in=5.671875 val=1.396281
    (addr==471) ? 23429658 :  //   in=5.679688 val=1.396517
    (addr==472) ? 23433594 :  //   in=5.687500 val=1.396751
    (addr==473) ? 23437519 :  //   in=5.695312 val=1.396985
    (addr==474) ? 23441434 :  //   in=5.703125 val=1.397218
    (addr==475) ? 23445339 :  //   in=5.710938 val=1.397451
    (addr==476) ? 23449233 :  //   in=5.718750 val=1.397683
    (addr==477) ? 23453116 :  //   in=5.726562 val=1.397915
    (addr==478) ? 23456990 :  //   in=5.734375 val=1.398146
    (addr==479) ? 23460853 :  //   in=5.742188 val=1.398376
    (addr==480) ? 23464706 :  //   in=5.750000 val=1.398606
    (addr==481) ? 23468549 :  //   in=5.757812 val=1.398835
    (addr==482) ? 23472382 :  //   in=5.765625 val=1.399063
    (addr==483) ? 23476205 :  //   in=5.773438 val=1.399291
    (addr==484) ? 23480017 :  //   in=5.781250 val=1.399518
    (addr==485) ? 23483820 :  //   in=5.789062 val=1.399745
    (addr==486) ? 23487613 :  //   in=5.796875 val=1.399971
    (addr==487) ? 23491396 :  //   in=5.804688 val=1.400196
    (addr==488) ? 23495169 :  //   in=5.812500 val=1.400421
    (addr==489) ? 23498932 :  //   in=5.820312 val=1.400646
    (addr==490) ? 23502685 :  //   in=5.828125 val=1.400869
    (addr==491) ? 23506429 :  //   in=5.835938 val=1.401092
    (addr==492) ? 23510163 :  //   in=5.843750 val=1.401315
    (addr==493) ? 23513887 :  //   in=5.851562 val=1.401537
    (addr==494) ? 23517601 :  //   in=5.859375 val=1.401758
    (addr==495) ? 23521306 :  //   in=5.867188 val=1.401979
    (addr==496) ? 23525001 :  //   in=5.875000 val=1.402199
    (addr==497) ? 23528687 :  //   in=5.882812 val=1.402419
    (addr==498) ? 23532364 :  //   in=5.890625 val=1.402638
    (addr==499) ? 23536030 :  //   in=5.898438 val=1.402857
    (addr==500) ? 23539688 :  //   in=5.906250 val=1.403075
    (addr==501) ? 23543336 :  //   in=5.914062 val=1.403292
    (addr==502) ? 23546974 :  //   in=5.921875 val=1.403509
    (addr==503) ? 23550604 :  //   in=5.929688 val=1.403725
    (addr==504) ? 23554224 :  //   in=5.937500 val=1.403941
    (addr==505) ? 23557834 :  //   in=5.945312 val=1.404156
    (addr==506) ? 23561436 :  //   in=5.953125 val=1.404371
    (addr==507) ? 23565028 :  //   in=5.960938 val=1.404585
    (addr==508) ? 23568612 :  //   in=5.968750 val=1.404799
    (addr==509) ? 23572186 :  //   in=5.976562 val=1.405012
    (addr==510) ? 23575751 :  //   in=5.984375 val=1.405224
    (addr==511) ? 23579307 :  //   in=5.992188 val=1.405436
    (addr==512) ? 23582854 :  //   in=6.000000 val=1.405648
    (addr==513) ? 23586392 :  //   in=6.007812 val=1.405859
    (addr==514) ? 23589921 :  //   in=6.015625 val=1.406069
    (addr==515) ? 23593441 :  //   in=6.023438 val=1.406279
    (addr==516) ? 23596952 :  //   in=6.031250 val=1.406488
    (addr==517) ? 23600455 :  //   in=6.039062 val=1.406697
    (addr==518) ? 23603948 :  //   in=6.046875 val=1.406905
    (addr==519) ? 23607433 :  //   in=6.054688 val=1.407113
    (addr==520) ? 23610909 :  //   in=6.062500 val=1.407320
    (addr==521) ? 23614377 :  //   in=6.070312 val=1.407527
    (addr==522) ? 23617835 :  //   in=6.078125 val=1.407733
    (addr==523) ? 23621285 :  //   in=6.085938 val=1.407938
    (addr==524) ? 23624727 :  //   in=6.093750 val=1.408143
    (addr==525) ? 23628160 :  //   in=6.101562 val=1.408348
    (addr==526) ? 23631584 :  //   in=6.109375 val=1.408552
    (addr==527) ? 23635000 :  //   in=6.117188 val=1.408756
    (addr==528) ? 23638407 :  //   in=6.125000 val=1.408959
    (addr==529) ? 23641806 :  //   in=6.132812 val=1.409161
    (addr==530) ? 23645197 :  //   in=6.140625 val=1.409364
    (addr==531) ? 23648579 :  //   in=6.148438 val=1.409565
    (addr==532) ? 23651952 :  //   in=6.156250 val=1.409766
    (addr==533) ? 23655318 :  //   in=6.164062 val=1.409967
    (addr==534) ? 23658675 :  //   in=6.171875 val=1.410167
    (addr==535) ? 23662023 :  //   in=6.179688 val=1.410367
    (addr==536) ? 23665364 :  //   in=6.187500 val=1.410566
    (addr==537) ? 23668696 :  //   in=6.195312 val=1.410764
    (addr==538) ? 23672020 :  //   in=6.203125 val=1.410962
    (addr==539) ? 23675336 :  //   in=6.210938 val=1.411160
    (addr==540) ? 23678644 :  //   in=6.218750 val=1.411357
    (addr==541) ? 23681944 :  //   in=6.226562 val=1.411554
    (addr==542) ? 23685236 :  //   in=6.234375 val=1.411750
    (addr==543) ? 23688519 :  //   in=6.242188 val=1.411946
    (addr==544) ? 23691795 :  //   in=6.250000 val=1.412141
    (addr==545) ? 23695063 :  //   in=6.257812 val=1.412336
    (addr==546) ? 23698323 :  //   in=6.265625 val=1.412530
    (addr==547) ? 23701574 :  //   in=6.273438 val=1.412724
    (addr==548) ? 23704818 :  //   in=6.281250 val=1.412917
    (addr==549) ? 23708055 :  //   in=6.289062 val=1.413110
    (addr==550) ? 23711283 :  //   in=6.296875 val=1.413303
    (addr==551) ? 23714503 :  //   in=6.304688 val=1.413495
    (addr==552) ? 23717716 :  //   in=6.312500 val=1.413686
    (addr==553) ? 23720921 :  //   in=6.320312 val=1.413877
    (addr==554) ? 23724118 :  //   in=6.328125 val=1.414068
    (addr==555) ? 23727308 :  //   in=6.335938 val=1.414258
    (addr==556) ? 23730489 :  //   in=6.343750 val=1.414447
    (addr==557) ? 23733664 :  //   in=6.351562 val=1.414637
    (addr==558) ? 23736830 :  //   in=6.359375 val=1.414825
    (addr==559) ? 23739989 :  //   in=6.367188 val=1.415014
    (addr==560) ? 23743141 :  //   in=6.375000 val=1.415201
    (addr==561) ? 23746285 :  //   in=6.382812 val=1.415389
    (addr==562) ? 23749421 :  //   in=6.390625 val=1.415576
    (addr==563) ? 23752550 :  //   in=6.398438 val=1.415762
    (addr==564) ? 23755672 :  //   in=6.406250 val=1.415948
    (addr==565) ? 23758786 :  //   in=6.414062 val=1.416134
    (addr==566) ? 23761892 :  //   in=6.421875 val=1.416319
    (addr==567) ? 23764992 :  //   in=6.429688 val=1.416504
    (addr==568) ? 23768084 :  //   in=6.437500 val=1.416688
    (addr==569) ? 23771168 :  //   in=6.445312 val=1.416872
    (addr==570) ? 23774246 :  //   in=6.453125 val=1.417055
    (addr==571) ? 23777316 :  //   in=6.460938 val=1.417238
    (addr==572) ? 23780379 :  //   in=6.468750 val=1.417421
    (addr==573) ? 23783434 :  //   in=6.476562 val=1.417603
    (addr==574) ? 23786483 :  //   in=6.484375 val=1.417785
    (addr==575) ? 23789524 :  //   in=6.492188 val=1.417966
    (addr==576) ? 23792558 :  //   in=6.500000 val=1.418147
    (addr==577) ? 23795585 :  //   in=6.507812 val=1.418327
    (addr==578) ? 23798605 :  //   in=6.515625 val=1.418507
    (addr==579) ? 23801618 :  //   in=6.523438 val=1.418687
    (addr==580) ? 23804624 :  //   in=6.531250 val=1.418866
    (addr==581) ? 23807622 :  //   in=6.539062 val=1.419045
    (addr==582) ? 23810614 :  //   in=6.546875 val=1.419223
    (addr==583) ? 23813599 :  //   in=6.554688 val=1.419401
    (addr==584) ? 23816577 :  //   in=6.562500 val=1.419579
    (addr==585) ? 23819548 :  //   in=6.570312 val=1.419756
    (addr==586) ? 23822512 :  //   in=6.578125 val=1.419932
    (addr==587) ? 23825469 :  //   in=6.585938 val=1.420109
    (addr==588) ? 23828419 :  //   in=6.593750 val=1.420285
    (addr==589) ? 23831363 :  //   in=6.601562 val=1.420460
    (addr==590) ? 23834300 :  //   in=6.609375 val=1.420635
    (addr==591) ? 23837230 :  //   in=6.617188 val=1.420810
    (addr==592) ? 23840153 :  //   in=6.625000 val=1.420984
    (addr==593) ? 23843069 :  //   in=6.632812 val=1.421158
    (addr==594) ? 23845979 :  //   in=6.640625 val=1.421331
    (addr==595) ? 23848882 :  //   in=6.648438 val=1.421504
    (addr==596) ? 23851778 :  //   in=6.656250 val=1.421677
    (addr==597) ? 23854668 :  //   in=6.664062 val=1.421849
    (addr==598) ? 23857551 :  //   in=6.671875 val=1.422021
    (addr==599) ? 23860428 :  //   in=6.679688 val=1.422192
    (addr==600) ? 23863298 :  //   in=6.687500 val=1.422363
    (addr==601) ? 23866161 :  //   in=6.695312 val=1.422534
    (addr==602) ? 23869018 :  //   in=6.703125 val=1.422704
    (addr==603) ? 23871868 :  //   in=6.710938 val=1.422874
    (addr==604) ? 23874712 :  //   in=6.718750 val=1.423044
    (addr==605) ? 23877550 :  //   in=6.726562 val=1.423213
    (addr==606) ? 23880381 :  //   in=6.734375 val=1.423382
    (addr==607) ? 23883205 :  //   in=6.742188 val=1.423550
    (addr==608) ? 23886023 :  //   in=6.750000 val=1.423718
    (addr==609) ? 23888835 :  //   in=6.757812 val=1.423886
    (addr==610) ? 23891641 :  //   in=6.765625 val=1.424053
    (addr==611) ? 23894440 :  //   in=6.773438 val=1.424220
    (addr==612) ? 23897233 :  //   in=6.781250 val=1.424386
    (addr==613) ? 23900019 :  //   in=6.789062 val=1.424552
    (addr==614) ? 23902799 :  //   in=6.796875 val=1.424718
    (addr==615) ? 23905573 :  //   in=6.804688 val=1.424883
    (addr==616) ? 23908341 :  //   in=6.812500 val=1.425048
    (addr==617) ? 23911103 :  //   in=6.820312 val=1.425213
    (addr==618) ? 23913858 :  //   in=6.828125 val=1.425377
    (addr==619) ? 23916607 :  //   in=6.835938 val=1.425541
    (addr==620) ? 23919350 :  //   in=6.843750 val=1.425704
    (addr==621) ? 23922087 :  //   in=6.851562 val=1.425868
    (addr==622) ? 23924818 :  //   in=6.859375 val=1.426030
    (addr==623) ? 23927543 :  //   in=6.867188 val=1.426193
    (addr==624) ? 23930261 :  //   in=6.875000 val=1.426355
    (addr==625) ? 23932974 :  //   in=6.882812 val=1.426516
    (addr==626) ? 23935680 :  //   in=6.890625 val=1.426678
    (addr==627) ? 23938381 :  //   in=6.898438 val=1.426839
    (addr==628) ? 23941076 :  //   in=6.906250 val=1.426999
    (addr==629) ? 23943764 :  //   in=6.914062 val=1.427160
    (addr==630) ? 23946447 :  //   in=6.921875 val=1.427319
    (addr==631) ? 23949124 :  //   in=6.929688 val=1.427479
    (addr==632) ? 23951795 :  //   in=6.937500 val=1.427638
    (addr==633) ? 23954460 :  //   in=6.945312 val=1.427797
    (addr==634) ? 23957119 :  //   in=6.953125 val=1.427956
    (addr==635) ? 23959772 :  //   in=6.960938 val=1.428114
    (addr==636) ? 23962419 :  //   in=6.968750 val=1.428272
    (addr==637) ? 23965061 :  //   in=6.976562 val=1.428429
    (addr==638) ? 23967697 :  //   in=6.984375 val=1.428586
    (addr==639) ? 23970327 :  //   in=6.992188 val=1.428743
    (addr==640) ? 23972951 :  //   in=7.000000 val=1.428899
    (addr==641) ? 23975570 :  //   in=7.007812 val=1.429055
    (addr==642) ? 23978183 :  //   in=7.015625 val=1.429211
    (addr==643) ? 23980790 :  //   in=7.023438 val=1.429366
    (addr==644) ? 23983391 :  //   in=7.031250 val=1.429522
    (addr==645) ? 23985987 :  //   in=7.039062 val=1.429676
    (addr==646) ? 23988577 :  //   in=7.046875 val=1.429831
    (addr==647) ? 23991162 :  //   in=7.054688 val=1.429985
    (addr==648) ? 23993741 :  //   in=7.062500 val=1.430138
    (addr==649) ? 23996314 :  //   in=7.070312 val=1.430292
    (addr==650) ? 23998882 :  //   in=7.078125 val=1.430445
    (addr==651) ? 24001444 :  //   in=7.085938 val=1.430598
    (addr==652) ? 24004001 :  //   in=7.093750 val=1.430750
    (addr==653) ? 24006552 :  //   in=7.101562 val=1.430902
    (addr==654) ? 24009098 :  //   in=7.109375 val=1.431054
    (addr==655) ? 24011638 :  //   in=7.117188 val=1.431205
    (addr==656) ? 24014173 :  //   in=7.125000 val=1.431356
    (addr==657) ? 24016702 :  //   in=7.132812 val=1.431507
    (addr==658) ? 24019226 :  //   in=7.140625 val=1.431657
    (addr==659) ? 24021744 :  //   in=7.148438 val=1.431808
    (addr==660) ? 24024258 :  //   in=7.156250 val=1.431957
    (addr==661) ? 24026765 :  //   in=7.164062 val=1.432107
    (addr==662) ? 24029268 :  //   in=7.171875 val=1.432256
    (addr==663) ? 24031765 :  //   in=7.179688 val=1.432405
    (addr==664) ? 24034256 :  //   in=7.187500 val=1.432553
    (addr==665) ? 24036743 :  //   in=7.195312 val=1.432702
    (addr==666) ? 24039224 :  //   in=7.203125 val=1.432849
    (addr==667) ? 24041699 :  //   in=7.210938 val=1.432997
    (addr==668) ? 24044170 :  //   in=7.218750 val=1.433144
    (addr==669) ? 24046635 :  //   in=7.226562 val=1.433291
    (addr==670) ? 24049095 :  //   in=7.234375 val=1.433438
    (addr==671) ? 24051550 :  //   in=7.242188 val=1.433584
    (addr==672) ? 24054000 :  //   in=7.250000 val=1.433730
    (addr==673) ? 24056444 :  //   in=7.257812 val=1.433876
    (addr==674) ? 24058884 :  //   in=7.265625 val=1.434021
    (addr==675) ? 24061318 :  //   in=7.273438 val=1.434166
    (addr==676) ? 24063747 :  //   in=7.281250 val=1.434311
    (addr==677) ? 24066171 :  //   in=7.289062 val=1.434456
    (addr==678) ? 24068590 :  //   in=7.296875 val=1.434600
    (addr==679) ? 24071004 :  //   in=7.304688 val=1.434744
    (addr==680) ? 24073412 :  //   in=7.312500 val=1.434887
    (addr==681) ? 24075816 :  //   in=7.320312 val=1.435030
    (addr==682) ? 24078215 :  //   in=7.328125 val=1.435173
    (addr==683) ? 24080608 :  //   in=7.335938 val=1.435316
    (addr==684) ? 24082997 :  //   in=7.343750 val=1.435459
    (addr==685) ? 24085381 :  //   in=7.351562 val=1.435601
    (addr==686) ? 24087759 :  //   in=7.359375 val=1.435742
    (addr==687) ? 24090133 :  //   in=7.367188 val=1.435884
    (addr==688) ? 24092502 :  //   in=7.375000 val=1.436025
    (addr==689) ? 24094866 :  //   in=7.382812 val=1.436166
    (addr==690) ? 24097225 :  //   in=7.390625 val=1.436307
    (addr==691) ? 24099579 :  //   in=7.398438 val=1.436447
    (addr==692) ? 24101928 :  //   in=7.406250 val=1.436587
    (addr==693) ? 24104272 :  //   in=7.414062 val=1.436727
    (addr==694) ? 24106612 :  //   in=7.421875 val=1.436866
    (addr==695) ? 24108946 :  //   in=7.429688 val=1.437005
    (addr==696) ? 24111276 :  //   in=7.437500 val=1.437144
    (addr==697) ? 24113601 :  //   in=7.445312 val=1.437283
    (addr==698) ? 24115921 :  //   in=7.453125 val=1.437421
    (addr==699) ? 24118237 :  //   in=7.460938 val=1.437559
    (addr==700) ? 24120548 :  //   in=7.468750 val=1.437697
    (addr==701) ? 24122854 :  //   in=7.476562 val=1.437834
    (addr==702) ? 24125155 :  //   in=7.484375 val=1.437971
    (addr==703) ? 24127451 :  //   in=7.492188 val=1.438108
    (addr==704) ? 24129743 :  //   in=7.500000 val=1.438245
    (addr==705) ? 24132030 :  //   in=7.507812 val=1.438381
    (addr==706) ? 24134313 :  //   in=7.515625 val=1.438517
    (addr==707) ? 24136590 :  //   in=7.523438 val=1.438653
    (addr==708) ? 24138864 :  //   in=7.531250 val=1.438788
    (addr==709) ? 24141132 :  //   in=7.539062 val=1.438924
    (addr==710) ? 24143396 :  //   in=7.546875 val=1.439059
    (addr==711) ? 24145655 :  //   in=7.554688 val=1.439193
    (addr==712) ? 24147910 :  //   in=7.562500 val=1.439328
    (addr==713) ? 24150160 :  //   in=7.570312 val=1.439462
    (addr==714) ? 24152406 :  //   in=7.578125 val=1.439596
    (addr==715) ? 24154647 :  //   in=7.585938 val=1.439729
    (addr==716) ? 24156883 :  //   in=7.593750 val=1.439862
    (addr==717) ? 24159115 :  //   in=7.601562 val=1.439996
    (addr==718) ? 24161343 :  //   in=7.609375 val=1.440128
    (addr==719) ? 24163566 :  //   in=7.617188 val=1.440261
    (addr==720) ? 24165784 :  //   in=7.625000 val=1.440393
    (addr==721) ? 24167998 :  //   in=7.632812 val=1.440525
    (addr==722) ? 24170208 :  //   in=7.640625 val=1.440657
    (addr==723) ? 24172413 :  //   in=7.648438 val=1.440788
    (addr==724) ? 24174614 :  //   in=7.656250 val=1.440919
    (addr==725) ? 24176810 :  //   in=7.664062 val=1.441050
    (addr==726) ? 24179002 :  //   in=7.671875 val=1.441181
    (addr==727) ? 24181190 :  //   in=7.679688 val=1.441311
    (addr==728) ? 24183373 :  //   in=7.687500 val=1.441441
    (addr==729) ? 24185552 :  //   in=7.695312 val=1.441571
    (addr==730) ? 24187726 :  //   in=7.703125 val=1.441701
    (addr==731) ? 24189896 :  //   in=7.710938 val=1.441830
    (addr==732) ? 24192062 :  //   in=7.718750 val=1.441959
    (addr==733) ? 24194223 :  //   in=7.726562 val=1.442088
    (addr==734) ? 24196381 :  //   in=7.734375 val=1.442217
    (addr==735) ? 24198534 :  //   in=7.742188 val=1.442345
    (addr==736) ? 24200682 :  //   in=7.750000 val=1.442473
    (addr==737) ? 24202827 :  //   in=7.757812 val=1.442601
    (addr==738) ? 24204967 :  //   in=7.765625 val=1.442728
    (addr==739) ? 24207103 :  //   in=7.773438 val=1.442856
    (addr==740) ? 24209234 :  //   in=7.781250 val=1.442983
    (addr==741) ? 24211362 :  //   in=7.789062 val=1.443110
    (addr==742) ? 24213485 :  //   in=7.796875 val=1.443236
    (addr==743) ? 24215604 :  //   in=7.804688 val=1.443363
    (addr==744) ? 24217719 :  //   in=7.812500 val=1.443489
    (addr==745) ? 24219830 :  //   in=7.820312 val=1.443614
    (addr==746) ? 24221937 :  //   in=7.828125 val=1.443740
    (addr==747) ? 24224039 :  //   in=7.835938 val=1.443865
    (addr==748) ? 24226138 :  //   in=7.843750 val=1.443990
    (addr==749) ? 24228232 :  //   in=7.851562 val=1.444115
    (addr==750) ? 24230322 :  //   in=7.859375 val=1.444240
    (addr==751) ? 24232408 :  //   in=7.867188 val=1.444364
    (addr==752) ? 24234490 :  //   in=7.875000 val=1.444488
    (addr==753) ? 24236568 :  //   in=7.882812 val=1.444612
    (addr==754) ? 24238642 :  //   in=7.890625 val=1.444736
    (addr==755) ? 24240712 :  //   in=7.898438 val=1.444859
    (addr==756) ? 24242778 :  //   in=7.906250 val=1.444982
    (addr==757) ? 24244840 :  //   in=7.914062 val=1.445105
    (addr==758) ? 24246897 :  //   in=7.921875 val=1.445228
    (addr==759) ? 24248951 :  //   in=7.929688 val=1.445350
    (addr==760) ? 24251001 :  //   in=7.937500 val=1.445472
    (addr==761) ? 24253047 :  //   in=7.945312 val=1.445594
    (addr==762) ? 24255089 :  //   in=7.953125 val=1.445716
    (addr==763) ? 24257127 :  //   in=7.960938 val=1.445837
    (addr==764) ? 24259161 :  //   in=7.968750 val=1.445959
    (addr==765) ? 24261191 :  //   in=7.976562 val=1.446080
    (addr==766) ? 24263217 :  //   in=7.984375 val=1.446200
    (addr==767) ? 24265240 :  //   in=7.992188 val=1.446321
    (addr==768) ? 24267258 :  //   in=8.000000 val=1.446441
    (addr==769) ? 24269273 :  //   in=8.007812 val=1.446561
    (addr==770) ? 24271283 :  //   in=8.015625 val=1.446681
    (addr==771) ? 24273290 :  //   in=8.023438 val=1.446801
    (addr==772) ? 24275293 :  //   in=8.031250 val=1.446920
    (addr==773) ? 24277292 :  //   in=8.039062 val=1.447039
    (addr==774) ? 24279288 :  //   in=8.046875 val=1.447158
    (addr==775) ? 24281279 :  //   in=8.054688 val=1.447277
    (addr==776) ? 24283267 :  //   in=8.062500 val=1.447396
    (addr==777) ? 24285251 :  //   in=8.070312 val=1.447514
    (addr==778) ? 24287231 :  //   in=8.078125 val=1.447632
    (addr==779) ? 24289207 :  //   in=8.085938 val=1.447750
    (addr==780) ? 24291180 :  //   in=8.093750 val=1.447867
    (addr==781) ? 24293149 :  //   in=8.101562 val=1.447985
    (addr==782) ? 24295114 :  //   in=8.109375 val=1.448102
    (addr==783) ? 24297075 :  //   in=8.117188 val=1.448219
    (addr==784) ? 24299033 :  //   in=8.125000 val=1.448335
    (addr==785) ? 24300987 :  //   in=8.132812 val=1.448452
    (addr==786) ? 24302937 :  //   in=8.140625 val=1.448568
    (addr==787) ? 24304884 :  //   in=8.148438 val=1.448684
    (addr==788) ? 24306827 :  //   in=8.156250 val=1.448800
    (addr==789) ? 24308766 :  //   in=8.164062 val=1.448915
    (addr==790) ? 24310702 :  //   in=8.171875 val=1.449031
    (addr==791) ? 24312634 :  //   in=8.179688 val=1.449146
    (addr==792) ? 24314562 :  //   in=8.187500 val=1.449261
    (addr==793) ? 24316487 :  //   in=8.195312 val=1.449376
    (addr==794) ? 24318408 :  //   in=8.203125 val=1.449490
    (addr==795) ? 24320326 :  //   in=8.210938 val=1.449604
    (addr==796) ? 24322239 :  //   in=8.218750 val=1.449718
    (addr==797) ? 24324150 :  //   in=8.226562 val=1.449832
    (addr==798) ? 24326057 :  //   in=8.234375 val=1.449946
    (addr==799) ? 24327960 :  //   in=8.242188 val=1.450059
    (addr==800) ? 24329859 :  //   in=8.250000 val=1.450173
    (addr==801) ? 24331756 :  //   in=8.257812 val=1.450286
    (addr==802) ? 24333648 :  //   in=8.265625 val=1.450398
    (addr==803) ? 24335537 :  //   in=8.273438 val=1.450511
    (addr==804) ? 24337423 :  //   in=8.281250 val=1.450623
    (addr==805) ? 24339305 :  //   in=8.289062 val=1.450736
    (addr==806) ? 24341183 :  //   in=8.296875 val=1.450848
    (addr==807) ? 24343058 :  //   in=8.304688 val=1.450959
    (addr==808) ? 24344930 :  //   in=8.312500 val=1.451071
    (addr==809) ? 24346798 :  //   in=8.320312 val=1.451182
    (addr==810) ? 24348663 :  //   in=8.328125 val=1.451293
    (addr==811) ? 24350524 :  //   in=8.335938 val=1.451404
    (addr==812) ? 24352382 :  //   in=8.343750 val=1.451515
    (addr==813) ? 24354236 :  //   in=8.351562 val=1.451626
    (addr==814) ? 24356087 :  //   in=8.359375 val=1.451736
    (addr==815) ? 24357935 :  //   in=8.367188 val=1.451846
    (addr==816) ? 24359779 :  //   in=8.375000 val=1.451956
    (addr==817) ? 24361619 :  //   in=8.382812 val=1.452066
    (addr==818) ? 24363457 :  //   in=8.390625 val=1.452175
    (addr==819) ? 24365291 :  //   in=8.398438 val=1.452285
    (addr==820) ? 24367121 :  //   in=8.406250 val=1.452394
    (addr==821) ? 24368949 :  //   in=8.414062 val=1.452503
    (addr==822) ? 24370773 :  //   in=8.421875 val=1.452611
    (addr==823) ? 24372593 :  //   in=8.429688 val=1.452720
    (addr==824) ? 24374410 :  //   in=8.437500 val=1.452828
    (addr==825) ? 24376224 :  //   in=8.445312 val=1.452936
    (addr==826) ? 24378035 :  //   in=8.453125 val=1.453044
    (addr==827) ? 24379842 :  //   in=8.460938 val=1.453152
    (addr==828) ? 24381646 :  //   in=8.468750 val=1.453259
    (addr==829) ? 24383447 :  //   in=8.476562 val=1.453367
    (addr==830) ? 24385245 :  //   in=8.484375 val=1.453474
    (addr==831) ? 24387039 :  //   in=8.492188 val=1.453581
    (addr==832) ? 24388830 :  //   in=8.500000 val=1.453688
    (addr==833) ? 24390618 :  //   in=8.507812 val=1.453794
    (addr==834) ? 24392402 :  //   in=8.515625 val=1.453901
    (addr==835) ? 24394184 :  //   in=8.523438 val=1.454007
    (addr==836) ? 24395962 :  //   in=8.531250 val=1.454113
    (addr==837) ? 24397737 :  //   in=8.539062 val=1.454218
    (addr==838) ? 24399508 :  //   in=8.546875 val=1.454324
    (addr==839) ? 24401277 :  //   in=8.554688 val=1.454429
    (addr==840) ? 24403042 :  //   in=8.562500 val=1.454535
    (addr==841) ? 24404804 :  //   in=8.570312 val=1.454640
    (addr==842) ? 24406563 :  //   in=8.578125 val=1.454745
    (addr==843) ? 24408319 :  //   in=8.585938 val=1.454849
    (addr==844) ? 24410072 :  //   in=8.593750 val=1.454954
    (addr==845) ? 24411821 :  //   in=8.601562 val=1.455058
    (addr==846) ? 24413567 :  //   in=8.609375 val=1.455162
    (addr==847) ? 24415311 :  //   in=8.617188 val=1.455266
    (addr==848) ? 24417051 :  //   in=8.625000 val=1.455370
    (addr==849) ? 24418788 :  //   in=8.632812 val=1.455473
    (addr==850) ? 24420522 :  //   in=8.640625 val=1.455577
    (addr==851) ? 24422253 :  //   in=8.648438 val=1.455680
    (addr==852) ? 24423980 :  //   in=8.656250 val=1.455783
    (addr==853) ? 24425705 :  //   in=8.664062 val=1.455885
    (addr==854) ? 24427427 :  //   in=8.671875 val=1.455988
    (addr==855) ? 24429145 :  //   in=8.679688 val=1.456091
    (addr==856) ? 24430861 :  //   in=8.687500 val=1.456193
    (addr==857) ? 24432573 :  //   in=8.695312 val=1.456295
    (addr==858) ? 24434282 :  //   in=8.703125 val=1.456397
    (addr==859) ? 24435989 :  //   in=8.710938 val=1.456498
    (addr==860) ? 24437692 :  //   in=8.718750 val=1.456600
    (addr==861) ? 24439393 :  //   in=8.726562 val=1.456701
    (addr==862) ? 24441090 :  //   in=8.734375 val=1.456803
    (addr==863) ? 24442784 :  //   in=8.742188 val=1.456904
    (addr==864) ? 24444476 :  //   in=8.750000 val=1.457004
    (addr==865) ? 24446164 :  //   in=8.757812 val=1.457105
    (addr==866) ? 24447850 :  //   in=8.765625 val=1.457205
    (addr==867) ? 24449532 :  //   in=8.773438 val=1.457306
    (addr==868) ? 24451211 :  //   in=8.781250 val=1.457406
    (addr==869) ? 24452888 :  //   in=8.789062 val=1.457506
    (addr==870) ? 24454562 :  //   in=8.796875 val=1.457605
    (addr==871) ? 24456232 :  //   in=8.804688 val=1.457705
    (addr==872) ? 24457900 :  //   in=8.812500 val=1.457804
    (addr==873) ? 24459565 :  //   in=8.820312 val=1.457904
    (addr==874) ? 24461227 :  //   in=8.828125 val=1.458003
    (addr==875) ? 24462886 :  //   in=8.835938 val=1.458102
    (addr==876) ? 24464542 :  //   in=8.843750 val=1.458200
    (addr==877) ? 24466195 :  //   in=8.851562 val=1.458299
    (addr==878) ? 24467846 :  //   in=8.859375 val=1.458397
    (addr==879) ? 24469493 :  //   in=8.867188 val=1.458495
    (addr==880) ? 24471138 :  //   in=8.875000 val=1.458594
    (addr==881) ? 24472780 :  //   in=8.882812 val=1.458691
    (addr==882) ? 24474419 :  //   in=8.890625 val=1.458789
    (addr==883) ? 24476055 :  //   in=8.898438 val=1.458887
    (addr==884) ? 24477688 :  //   in=8.906250 val=1.458984
    (addr==885) ? 24479318 :  //   in=8.914062 val=1.459081
    (addr==886) ? 24480946 :  //   in=8.921875 val=1.459178
    (addr==887) ? 24482571 :  //   in=8.929688 val=1.459275
    (addr==888) ? 24484193 :  //   in=8.937500 val=1.459372
    (addr==889) ? 24485812 :  //   in=8.945312 val=1.459468
    (addr==890) ? 24487428 :  //   in=8.953125 val=1.459565
    (addr==891) ? 24489042 :  //   in=8.960938 val=1.459661
    (addr==892) ? 24490653 :  //   in=8.968750 val=1.459757
    (addr==893) ? 24492261 :  //   in=8.976562 val=1.459853
    (addr==894) ? 24493866 :  //   in=8.984375 val=1.459948
    (addr==895) ? 24495469 :  //   in=8.992188 val=1.460044
    (addr==896) ? 24497069 :  //   in=9.000000 val=1.460139
    (addr==897) ? 24498666 :  //   in=9.007812 val=1.460234
    (addr==898) ? 24500260 :  //   in=9.015625 val=1.460329
    (addr==899) ? 24501852 :  //   in=9.023438 val=1.460424
    (addr==900) ? 24503441 :  //   in=9.031250 val=1.460519
    (addr==901) ? 24505027 :  //   in=9.039062 val=1.460613
    (addr==902) ? 24506610 :  //   in=9.046875 val=1.460708
    (addr==903) ? 24508191 :  //   in=9.054688 val=1.460802
    (addr==904) ? 24509769 :  //   in=9.062500 val=1.460896
    (addr==905) ? 24511344 :  //   in=9.070312 val=1.460990
    (addr==906) ? 24512917 :  //   in=9.078125 val=1.461084
    (addr==907) ? 24514487 :  //   in=9.085938 val=1.461177
    (addr==908) ? 24516055 :  //   in=9.093750 val=1.461271
    (addr==909) ? 24517619 :  //   in=9.101562 val=1.461364
    (addr==910) ? 24519181 :  //   in=9.109375 val=1.461457
    (addr==911) ? 24520741 :  //   in=9.117188 val=1.461550
    (addr==912) ? 24522298 :  //   in=9.125000 val=1.461643
    (addr==913) ? 24523852 :  //   in=9.132812 val=1.461735
    (addr==914) ? 24525403 :  //   in=9.140625 val=1.461828
    (addr==915) ? 24526952 :  //   in=9.148438 val=1.461920
    (addr==916) ? 24528498 :  //   in=9.156250 val=1.462012
    (addr==917) ? 24530042 :  //   in=9.164062 val=1.462104
    (addr==918) ? 24531583 :  //   in=9.171875 val=1.462196
    (addr==919) ? 24533122 :  //   in=9.179688 val=1.462288
    (addr==920) ? 24534658 :  //   in=9.187500 val=1.462380
    (addr==921) ? 24536191 :  //   in=9.195312 val=1.462471
    (addr==922) ? 24537722 :  //   in=9.203125 val=1.462562
    (addr==923) ? 24539250 :  //   in=9.210938 val=1.462653
    (addr==924) ? 24540775 :  //   in=9.218750 val=1.462744
    (addr==925) ? 24542299 :  //   in=9.226562 val=1.462835
    (addr==926) ? 24543819 :  //   in=9.234375 val=1.462926
    (addr==927) ? 24545337 :  //   in=9.242188 val=1.463016
    (addr==928) ? 24546853 :  //   in=9.250000 val=1.463106
    (addr==929) ? 24548365 :  //   in=9.257812 val=1.463197
    (addr==930) ? 24549876 :  //   in=9.265625 val=1.463287
    (addr==931) ? 24551384 :  //   in=9.273438 val=1.463377
    (addr==932) ? 24552889 :  //   in=9.281250 val=1.463466
    (addr==933) ? 24554392 :  //   in=9.289062 val=1.463556
    (addr==934) ? 24555892 :  //   in=9.296875 val=1.463645
    (addr==935) ? 24557390 :  //   in=9.304688 val=1.463735
    (addr==936) ? 24558886 :  //   in=9.312500 val=1.463824
    (addr==937) ? 24560379 :  //   in=9.320312 val=1.463913
    (addr==938) ? 24561869 :  //   in=9.328125 val=1.464002
    (addr==939) ? 24563357 :  //   in=9.335938 val=1.464090
    (addr==940) ? 24564843 :  //   in=9.343750 val=1.464179
    (addr==941) ? 24566326 :  //   in=9.351562 val=1.464267
    (addr==942) ? 24567806 :  //   in=9.359375 val=1.464355
    (addr==943) ? 24569284 :  //   in=9.367188 val=1.464444
    (addr==944) ? 24570760 :  //   in=9.375000 val=1.464531
    (addr==945) ? 24572234 :  //   in=9.382812 val=1.464619
    (addr==946) ? 24573704 :  //   in=9.390625 val=1.464707
    (addr==947) ? 24575173 :  //   in=9.398438 val=1.464794
    (addr==948) ? 24576639 :  //   in=9.406250 val=1.464882
    (addr==949) ? 24578103 :  //   in=9.414062 val=1.464969
    (addr==950) ? 24579564 :  //   in=9.421875 val=1.465056
    (addr==951) ? 24581023 :  //   in=9.429688 val=1.465143
    (addr==952) ? 24582479 :  //   in=9.437500 val=1.465230
    (addr==953) ? 24583933 :  //   in=9.445312 val=1.465317
    (addr==954) ? 24585385 :  //   in=9.453125 val=1.465403
    (addr==955) ? 24586834 :  //   in=9.460938 val=1.465490
    (addr==956) ? 24588281 :  //   in=9.468750 val=1.465576
    (addr==957) ? 24589726 :  //   in=9.476562 val=1.465662
    (addr==958) ? 24591168 :  //   in=9.484375 val=1.465748
    (addr==959) ? 24592608 :  //   in=9.492188 val=1.465834
    (addr==960) ? 24594046 :  //   in=9.500000 val=1.465919
    (addr==961) ? 24595481 :  //   in=9.507812 val=1.466005
    (addr==962) ? 24596914 :  //   in=9.515625 val=1.466090
    (addr==963) ? 24598344 :  //   in=9.523438 val=1.466176
    (addr==964) ? 24599773 :  //   in=9.531250 val=1.466261
    (addr==965) ? 24601199 :  //   in=9.539062 val=1.466346
    (addr==966) ? 24602622 :  //   in=9.546875 val=1.466431
    (addr==967) ? 24604044 :  //   in=9.554688 val=1.466515
    (addr==968) ? 24605463 :  //   in=9.562500 val=1.466600
    (addr==969) ? 24606879 :  //   in=9.570312 val=1.466684
    (addr==970) ? 24608294 :  //   in=9.578125 val=1.466769
    (addr==971) ? 24609706 :  //   in=9.585938 val=1.466853
    (addr==972) ? 24611116 :  //   in=9.593750 val=1.466937
    (addr==973) ? 24612524 :  //   in=9.601562 val=1.467021
    (addr==974) ? 24613929 :  //   in=9.609375 val=1.467105
    (addr==975) ? 24615332 :  //   in=9.617188 val=1.467188
    (addr==976) ? 24616733 :  //   in=9.625000 val=1.467272
    (addr==977) ? 24618132 :  //   in=9.632812 val=1.467355
    (addr==978) ? 24619528 :  //   in=9.640625 val=1.467438
    (addr==979) ? 24620922 :  //   in=9.648438 val=1.467521
    (addr==980) ? 24622314 :  //   in=9.656250 val=1.467604
    (addr==981) ? 24623704 :  //   in=9.664062 val=1.467687
    (addr==982) ? 24625091 :  //   in=9.671875 val=1.467770
    (addr==983) ? 24626476 :  //   in=9.679688 val=1.467852
    (addr==984) ? 24627859 :  //   in=9.687500 val=1.467935
    (addr==985) ? 24629240 :  //   in=9.695312 val=1.468017
    (addr==986) ? 24630619 :  //   in=9.703125 val=1.468099
    (addr==987) ? 24631995 :  //   in=9.710938 val=1.468181
    (addr==988) ? 24633369 :  //   in=9.718750 val=1.468263
    (addr==989) ? 24634741 :  //   in=9.726562 val=1.468345
    (addr==990) ? 24636111 :  //   in=9.734375 val=1.468427
    (addr==991) ? 24637479 :  //   in=9.742188 val=1.468508
    (addr==992) ? 24638845 :  //   in=9.750000 val=1.468590
    (addr==993) ? 24640208 :  //   in=9.757812 val=1.468671
    (addr==994) ? 24641569 :  //   in=9.765625 val=1.468752
    (addr==995) ? 24642928 :  //   in=9.773438 val=1.468833
    (addr==996) ? 24644285 :  //   in=9.781250 val=1.468914
    (addr==997) ? 24645640 :  //   in=9.789062 val=1.468995
    (addr==998) ? 24646992 :  //   in=9.796875 val=1.469075
    (addr==999) ? 24648343 :  //   in=9.804688 val=1.469156
    (addr==1000) ? 24649691 :  //   in=9.812500 val=1.469236
    (addr==1001) ? 24651038 :  //   in=9.820312 val=1.469316
    (addr==1002) ? 24652382 :  //   in=9.828125 val=1.469396
    (addr==1003) ? 24653724 :  //   in=9.835938 val=1.469476
    (addr==1004) ? 24655064 :  //   in=9.843750 val=1.469556
    (addr==1005) ? 24656401 :  //   in=9.851562 val=1.469636
    (addr==1006) ? 24657737 :  //   in=9.859375 val=1.469716
    (addr==1007) ? 24659071 :  //   in=9.867188 val=1.469795
    (addr==1008) ? 24660402 :  //   in=9.875000 val=1.469875
    (addr==1009) ? 24661732 :  //   in=9.882812 val=1.469954
    (addr==1010) ? 24663059 :  //   in=9.890625 val=1.470033
    (addr==1011) ? 24664384 :  //   in=9.898438 val=1.470112
    (addr==1012) ? 24665707 :  //   in=9.906250 val=1.470191
    (addr==1013) ? 24667029 :  //   in=9.914062 val=1.470270
    (addr==1014) ? 24668348 :  //   in=9.921875 val=1.470348
    (addr==1015) ? 24669665 :  //   in=9.929688 val=1.470427
    (addr==1016) ? 24670980 :  //   in=9.937500 val=1.470505
    (addr==1017) ? 24672293 :  //   in=9.945312 val=1.470583
    (addr==1018) ? 24673603 :  //   in=9.953125 val=1.470661
    (addr==1019) ? 24674912 :  //   in=9.960938 val=1.470739
    (addr==1020) ? 24676219 :  //   in=9.968750 val=1.470817
    (addr==1021) ? 24677524 :  //   in=9.976562 val=1.470895
    (addr==1022) ? 24678827 :  //   in=9.984375 val=1.470973
    (addr==1023) ? 24680128 :  //   in=9.992188 val=1.471050
25'bx;
assign lastone = 24681426;
endmodule
