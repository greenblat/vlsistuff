`define RGF2_BASEADDR    'h0
`define ADDR_REGA                                                'h40000
`define ADDR_CONTROL0                                            'h40004
`define ADDR_STATUSA                                             'h40008
`define ADDR_REGB                                                'h4000c
`define ADDR_EXTERN                                              'h40010
`define ADDR_ETH0TMP0                                            'h40100
`define ADDR_ETH0TMP1                                            'h40104
`define ADDR_ETH0TMP2                                            'h40108
`define ADDR_ETH1TMP0                                            'h40200
`define ADDR_ETH1TMP1                                            'h40204
`define ADDR_ETH1TMP2                                            'h40208
`define ADDR_ETH2TMP0                                            'h40300
`define ADDR_ETH2TMP1                                            'h40304
`define ADDR_ETH2TMP2                                            'h40308
`define ADDR_ETH3TMP0                                            'h40400
`define ADDR_ETH3TMP1                                            'h40404
`define ADDR_ETH3TMP2                                            'h40408
`define ADDR_WIDER                                               'h4040c
`define ADDR_LONGER                                              'h4041c
`define ADDR_RONLY                                               'h4042c
`define ADDR_RONLY2                                              'h40430
`define ADDR_LDST_RAM                                            'h40800
