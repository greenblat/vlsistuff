`define FIR_RGF_BASEADDR    'h0
`define ADDR_ENABLE                                              'h0
`define ADDR_SCALEFACTOR                                         'h4
`define ADDR_COEFFS                                              'h8
`define ADDR_GOODS                                               'h28
`define ADDR_BADS                                                'h2c
