module sqrt_u48_6 ( input clk,input rst_n,input en,input vldin, input [47:0] ain, output reg [23:0] out,output reg vldout);
  // stages=6 places=[19, 14, 9, 4]
  // reg vld24;
  // always @(posedge clk) if (en) vld24 <= vldin;
  // reg [47:0] datain24;
  // always @(posedge clk) if (en) datain24 <= ain;
wire vld24 = vldin;
wire [47:0] datain24 = ain;
wire [47:0] Y24 = 0;
wire [47:0] YY24 = 0;
wire [47:0] Decra23 = (48'b1<<(2*23));
wire [47:0] Decrb23 = (Y24<<(23+1));
wire [47:0] Decr23 = Decra23+Decrb23;
wire [47:0] YY23_1 = YY24+Decr23;
wire [47:0] Base23 =  48'b1<<23;
wire smaller23 =  (YY23_1<=datain24);
wire [47:0] YY23 = smaller23 ? YY23_1 : YY24;
wire [23:0] Y23 = smaller23 ? Y24+Base23 : Y24;
wire [47:0] datain23 = datain24;
wire vld23 = vld24;
wire [47:0] Decra22 = (48'b1<<(2*22));
wire [47:0] Decrb22 = (Y23<<(22+1));
wire [47:0] Decr22 = Decra22+Decrb22;
wire [47:0] YY22_1 = YY23+Decr22;
wire [47:0] Base22 =  48'b1<<22;
wire smaller22 =  (YY22_1<=datain23);
wire [47:0] YY22 = smaller22 ? YY22_1 : YY23;
wire [23:0] Y22 = smaller22 ? Y23+Base22 : Y23;
wire [47:0] datain22 = datain23;
wire vld22 = vld23;
wire [47:0] Decra21 = (48'b1<<(2*21));
wire [47:0] Decrb21 = (Y22<<(21+1));
wire [47:0] Decr21 = Decra21+Decrb21;
wire [47:0] YY21_1 = YY22+Decr21;
wire [47:0] Base21 =  48'b1<<21;
wire smaller21 =  (YY21_1<=datain22);
wire [47:0] YY21 = smaller21 ? YY21_1 : YY22;
wire [23:0] Y21 = smaller21 ? Y22+Base21 : Y22;
wire [47:0] datain21 = datain22;
wire vld21 = vld22;
wire [47:0] Decra20 = (48'b1<<(2*20));
wire [47:0] Decrb20 = (Y21<<(20+1));
wire [47:0] Decr20 = Decra20+Decrb20;
wire [47:0] YY20_1 = YY21+Decr20;
wire [47:0] Base20 =  48'b1<<20;
wire smaller20 =  (YY20_1<=datain21);
wire [47:0] YY20 = smaller20 ? YY20_1 : YY21;
wire [23:0] Y20 = smaller20 ? Y21+Base20 : Y21;
wire [47:0] datain20 = datain21;
wire vld20 = vld21;
wire [47:0] Decra19 = (48'b1<<(2*19));
wire [47:0] Decrb19 = (Y20<<(19+1));
wire [47:0] Decr19 = Decra19+Decrb19;
wire [47:0] YY19_1 = YY20+Decr19;
wire [47:0] Base19 =  48'b1<<19;
wire smaller19 =  (YY19_1<=datain20);
wire [47:0] pre_YY19 = smaller19 ? YY19_1 : YY20;
wire [23:0] pre_Y19 = smaller19 ? Y20+Base19 : Y20;
reg [47:0] YY19;
always @(posedge clk) if (en) YY19 <= pre_YY19;
reg [47:0] Y19;
always @(posedge clk) if (en) Y19 <= pre_Y19;
reg [47:0] datain19;
always @(posedge clk) if (en) datain19 <= datain20;
reg vld19;
always @(posedge clk) if (en) vld19 <= vld20;
wire [47:0] Decra18 = (48'b1<<(2*18));
wire [47:0] Decrb18 = (Y19<<(18+1));
wire [47:0] Decr18 = Decra18+Decrb18;
wire [47:0] YY18_1 = YY19+Decr18;
wire [47:0] Base18 =  48'b1<<18;
wire smaller18 =  (YY18_1<=datain19);
wire [47:0] YY18 = smaller18 ? YY18_1 : YY19;
wire [23:0] Y18 = smaller18 ? Y19+Base18 : Y19;
wire [47:0] datain18 = datain19;
wire vld18 = vld19;
wire [47:0] Decra17 = (48'b1<<(2*17));
wire [47:0] Decrb17 = (Y18<<(17+1));
wire [47:0] Decr17 = Decra17+Decrb17;
wire [47:0] YY17_1 = YY18+Decr17;
wire [47:0] Base17 =  48'b1<<17;
wire smaller17 =  (YY17_1<=datain18);
wire [47:0] YY17 = smaller17 ? YY17_1 : YY18;
wire [23:0] Y17 = smaller17 ? Y18+Base17 : Y18;
wire [47:0] datain17 = datain18;
wire vld17 = vld18;
wire [47:0] Decra16 = (48'b1<<(2*16));
wire [47:0] Decrb16 = (Y17<<(16+1));
wire [47:0] Decr16 = Decra16+Decrb16;
wire [47:0] YY16_1 = YY17+Decr16;
wire [47:0] Base16 =  48'b1<<16;
wire smaller16 =  (YY16_1<=datain17);
wire [47:0] YY16 = smaller16 ? YY16_1 : YY17;
wire [23:0] Y16 = smaller16 ? Y17+Base16 : Y17;
wire [47:0] datain16 = datain17;
wire vld16 = vld17;
wire [47:0] Decra15 = (48'b1<<(2*15));
wire [47:0] Decrb15 = (Y16<<(15+1));
wire [47:0] Decr15 = Decra15+Decrb15;
wire [47:0] YY15_1 = YY16+Decr15;
wire [47:0] Base15 =  48'b1<<15;
wire smaller15 =  (YY15_1<=datain16);
wire [47:0] YY15 = smaller15 ? YY15_1 : YY16;
wire [23:0] Y15 = smaller15 ? Y16+Base15 : Y16;
wire [47:0] datain15 = datain16;
wire vld15 = vld16;
wire [47:0] Decra14 = (48'b1<<(2*14));
wire [47:0] Decrb14 = (Y15<<(14+1));
wire [47:0] Decr14 = Decra14+Decrb14;
wire [47:0] YY14_1 = YY15+Decr14;
wire [47:0] Base14 =  48'b1<<14;
wire smaller14 =  (YY14_1<=datain15);
wire [47:0] pre_YY14 = smaller14 ? YY14_1 : YY15;
wire [23:0] pre_Y14 = smaller14 ? Y15+Base14 : Y15;
reg [47:0] YY14;
always @(posedge clk) if (en) YY14 <= pre_YY14;
reg [47:0] Y14;
always @(posedge clk) if (en) Y14 <= pre_Y14;
reg [47:0] datain14;
always @(posedge clk) if (en) datain14 <= datain15;
reg vld14;
always @(posedge clk) if (en) vld14 <= vld15;
wire [47:0] Decra13 = (48'b1<<(2*13));
wire [47:0] Decrb13 = (Y14<<(13+1));
wire [47:0] Decr13 = Decra13+Decrb13;
wire [47:0] YY13_1 = YY14+Decr13;
wire [47:0] Base13 =  48'b1<<13;
wire smaller13 =  (YY13_1<=datain14);
wire [47:0] YY13 = smaller13 ? YY13_1 : YY14;
wire [23:0] Y13 = smaller13 ? Y14+Base13 : Y14;
wire [47:0] datain13 = datain14;
wire vld13 = vld14;
wire [47:0] Decra12 = (48'b1<<(2*12));
wire [47:0] Decrb12 = (Y13<<(12+1));
wire [47:0] Decr12 = Decra12+Decrb12;
wire [47:0] YY12_1 = YY13+Decr12;
wire [47:0] Base12 =  48'b1<<12;
wire smaller12 =  (YY12_1<=datain13);
wire [47:0] YY12 = smaller12 ? YY12_1 : YY13;
wire [23:0] Y12 = smaller12 ? Y13+Base12 : Y13;
wire [47:0] datain12 = datain13;
wire vld12 = vld13;
wire [47:0] Decra11 = (48'b1<<(2*11));
wire [47:0] Decrb11 = (Y12<<(11+1));
wire [47:0] Decr11 = Decra11+Decrb11;
wire [47:0] YY11_1 = YY12+Decr11;
wire [47:0] Base11 =  48'b1<<11;
wire smaller11 =  (YY11_1<=datain12);
wire [47:0] YY11 = smaller11 ? YY11_1 : YY12;
wire [23:0] Y11 = smaller11 ? Y12+Base11 : Y12;
wire [47:0] datain11 = datain12;
wire vld11 = vld12;
wire [47:0] Decra10 = (48'b1<<(2*10));
wire [47:0] Decrb10 = (Y11<<(10+1));
wire [47:0] Decr10 = Decra10+Decrb10;
wire [47:0] YY10_1 = YY11+Decr10;
wire [47:0] Base10 =  48'b1<<10;
wire smaller10 =  (YY10_1<=datain11);
wire [47:0] YY10 = smaller10 ? YY10_1 : YY11;
wire [23:0] Y10 = smaller10 ? Y11+Base10 : Y11;
wire [47:0] datain10 = datain11;
wire vld10 = vld11;
wire [47:0] Decra9 = (48'b1<<(2*9));
wire [47:0] Decrb9 = (Y10<<(9+1));
wire [47:0] Decr9 = Decra9+Decrb9;
wire [47:0] YY9_1 = YY10+Decr9;
wire [47:0] Base9 =  48'b1<<9;
wire smaller9 =  (YY9_1<=datain10);
wire [47:0] pre_YY9 = smaller9 ? YY9_1 : YY10;
wire [23:0] pre_Y9 = smaller9 ? Y10+Base9 : Y10;
reg [47:0] YY9;
always @(posedge clk) if (en) YY9 <= pre_YY9;
reg [47:0] Y9;
always @(posedge clk) if (en) Y9 <= pre_Y9;
reg [47:0] datain9;
always @(posedge clk) if (en) datain9 <= datain10;
reg vld9;
always @(posedge clk) if (en) vld9 <= vld10;
wire [47:0] Decra8 = (48'b1<<(2*8));
wire [47:0] Decrb8 = (Y9<<(8+1));
wire [47:0] Decr8 = Decra8+Decrb8;
wire [47:0] YY8_1 = YY9+Decr8;
wire [47:0] Base8 =  48'b1<<8;
wire smaller8 =  (YY8_1<=datain9);
wire [47:0] YY8 = smaller8 ? YY8_1 : YY9;
wire [23:0] Y8 = smaller8 ? Y9+Base8 : Y9;
wire [47:0] datain8 = datain9;
wire vld8 = vld9;
wire [47:0] Decra7 = (48'b1<<(2*7));
wire [47:0] Decrb7 = (Y8<<(7+1));
wire [47:0] Decr7 = Decra7+Decrb7;
wire [47:0] YY7_1 = YY8+Decr7;
wire [47:0] Base7 =  48'b1<<7;
wire smaller7 =  (YY7_1<=datain8);
wire [47:0] YY7 = smaller7 ? YY7_1 : YY8;
wire [23:0] Y7 = smaller7 ? Y8+Base7 : Y8;
wire [47:0] datain7 = datain8;
wire vld7 = vld8;
wire [47:0] Decra6 = (48'b1<<(2*6));
wire [47:0] Decrb6 = (Y7<<(6+1));
wire [47:0] Decr6 = Decra6+Decrb6;
wire [47:0] YY6_1 = YY7+Decr6;
wire [47:0] Base6 =  48'b1<<6;
wire smaller6 =  (YY6_1<=datain7);
wire [47:0] YY6 = smaller6 ? YY6_1 : YY7;
wire [23:0] Y6 = smaller6 ? Y7+Base6 : Y7;
wire [47:0] datain6 = datain7;
wire vld6 = vld7;
wire [47:0] Decra5 = (48'b1<<(2*5));
wire [47:0] Decrb5 = (Y6<<(5+1));
wire [47:0] Decr5 = Decra5+Decrb5;
wire [47:0] YY5_1 = YY6+Decr5;
wire [47:0] Base5 =  48'b1<<5;
wire smaller5 =  (YY5_1<=datain6);
wire [47:0] YY5 = smaller5 ? YY5_1 : YY6;
wire [23:0] Y5 = smaller5 ? Y6+Base5 : Y6;
wire [47:0] datain5 = datain6;
wire vld5 = vld6;
wire [47:0] Decra4 = (48'b1<<(2*4));
wire [47:0] Decrb4 = (Y5<<(4+1));
wire [47:0] Decr4 = Decra4+Decrb4;
wire [47:0] YY4_1 = YY5+Decr4;
wire [47:0] Base4 =  48'b1<<4;
wire smaller4 =  (YY4_1<=datain5);
wire [47:0] pre_YY4 = smaller4 ? YY4_1 : YY5;
wire [23:0] pre_Y4 = smaller4 ? Y5+Base4 : Y5;
reg [47:0] YY4;
always @(posedge clk) if (en) YY4 <= pre_YY4;
reg [47:0] Y4;
always @(posedge clk) if (en) Y4 <= pre_Y4;
reg [47:0] datain4;
always @(posedge clk) if (en) datain4 <= datain5;
reg vld4;
always @(posedge clk) if (en) vld4 <= vld5;
wire [47:0] Decra3 = (48'b1<<(2*3));
wire [47:0] Decrb3 = (Y4<<(3+1));
wire [47:0] Decr3 = Decra3+Decrb3;
wire [47:0] YY3_1 = YY4+Decr3;
wire [47:0] Base3 =  48'b1<<3;
wire smaller3 =  (YY3_1<=datain4);
wire [47:0] YY3 = smaller3 ? YY3_1 : YY4;
wire [23:0] Y3 = smaller3 ? Y4+Base3 : Y4;
wire [47:0] datain3 = datain4;
wire vld3 = vld4;
wire [47:0] Decra2 = (48'b1<<(2*2));
wire [47:0] Decrb2 = (Y3<<(2+1));
wire [47:0] Decr2 = Decra2+Decrb2;
wire [47:0] YY2_1 = YY3+Decr2;
wire [47:0] Base2 =  48'b1<<2;
wire smaller2 =  (YY2_1<=datain3);
wire [47:0] YY2 = smaller2 ? YY2_1 : YY3;
wire [23:0] Y2 = smaller2 ? Y3+Base2 : Y3;
wire [47:0] datain2 = datain3;
wire vld2 = vld3;
wire [47:0] Decra1 = (48'b1<<(2*1));
wire [47:0] Decrb1 = (Y2<<(1+1));
wire [47:0] Decr1 = Decra1+Decrb1;
wire [47:0] YY1_1 = YY2+Decr1;
wire [47:0] Base1 =  48'b1<<1;
wire smaller1 =  (YY1_1<=datain2);
wire [47:0] YY1 = smaller1 ? YY1_1 : YY2;
wire [23:0] Y1 = smaller1 ? Y2+Base1 : Y2;
wire [47:0] datain1 = datain2;
wire vld1 = vld2;
wire [47:0] Decra0 = (48'b1<<(2*0));
wire [47:0] Decrb0 = (Y1<<(0+1));
wire [47:0] Decr0 = Decra0+Decrb0;
wire [47:0] YY0_1 = YY1+Decr0;
wire [47:0] Base0 =  48'b1<<0;
wire smaller0 =  (YY0_1<=datain1);
wire [47:0] YY0 = smaller0 ? YY0_1 : YY1;
wire [23:0] Y0 = smaller0 ? Y1+Base0 : Y1;
wire [47:0] datain0 = datain1;
wire vld0 = vld1;
always @(posedge clk) if (en) out <= Y0;
always @(posedge clk) if (en) vldout <= vld0;
endmodule
