module example0(
    input  clk
    ,input [7:0] inx
    ,output reg [7:0] outx
    ,input  rst_n
);
endmodule

