module asin_table(input [9:0] addr,output [24:0] result);
assign result = 
    (addr==0) ? 0 :
    (addr==1) ? 16384 :
    (addr==2) ? 32768 :
    (addr==3) ? 49152 :
    (addr==4) ? 65536 :
    (addr==5) ? 81920 :
    (addr==6) ? 98304 :
    (addr==7) ? 114688 :
    (addr==8) ? 131073 :
    (addr==9) ? 147457 :
    (addr==10) ? 163842 :
    (addr==11) ? 180227 :
    (addr==12) ? 196612 :
    (addr==13) ? 212997 :
    (addr==14) ? 229383 :
    (addr==15) ? 245768 :
    (addr==16) ? 262154 :
    (addr==17) ? 278540 :
    (addr==18) ? 294927 :
    (addr==19) ? 311313 :
    (addr==20) ? 327700 :
    (addr==21) ? 344088 :
    (addr==22) ? 360475 :
    (addr==23) ? 376863 :
    (addr==24) ? 393252 :
    (addr==25) ? 409640 :
    (addr==26) ? 426029 :
    (addr==27) ? 442419 :
    (addr==28) ? 458809 :
    (addr==29) ? 475199 :
    (addr==30) ? 491590 :
    (addr==31) ? 507981 :
    (addr==32) ? 524373 :
    (addr==33) ? 540765 :
    (addr==34) ? 557158 :
    (addr==35) ? 573551 :
    (addr==36) ? 589945 :
    (addr==37) ? 606339 :
    (addr==38) ? 622734 :
    (addr==39) ? 639130 :
    (addr==40) ? 655526 :
    (addr==41) ? 671923 :
    (addr==42) ? 688321 :
    (addr==43) ? 704719 :
    (addr==44) ? 721118 :
    (addr==45) ? 737517 :
    (addr==46) ? 753917 :
    (addr==47) ? 770318 :
    (addr==48) ? 786720 :
    (addr==49) ? 803122 :
    (addr==50) ? 819525 :
    (addr==51) ? 835929 :
    (addr==52) ? 852334 :
    (addr==53) ? 868740 :
    (addr==54) ? 885146 :
    (addr==55) ? 901553 :
    (addr==56) ? 917961 :
    (addr==57) ? 934370 :
    (addr==58) ? 950780 :
    (addr==59) ? 967191 :
    (addr==60) ? 983603 :
    (addr==61) ? 1000016 :
    (addr==62) ? 1016429 :
    (addr==63) ? 1032844 :
    (addr==64) ? 1049259 :
    (addr==65) ? 1065676 :
    (addr==66) ? 1082094 :
    (addr==67) ? 1098512 :
    (addr==68) ? 1114932 :
    (addr==69) ? 1131353 :
    (addr==70) ? 1147775 :
    (addr==71) ? 1164198 :
    (addr==72) ? 1180622 :
    (addr==73) ? 1197047 :
    (addr==74) ? 1213473 :
    (addr==75) ? 1229901 :
    (addr==76) ? 1246330 :
    (addr==77) ? 1262759 :
    (addr==78) ? 1279191 :
    (addr==79) ? 1295623 :
    (addr==80) ? 1312057 :
    (addr==81) ? 1328491 :
    (addr==82) ? 1344928 :
    (addr==83) ? 1361365 :
    (addr==84) ? 1377804 :
    (addr==85) ? 1394244 :
    (addr==86) ? 1410685 :
    (addr==87) ? 1427128 :
    (addr==88) ? 1443572 :
    (addr==89) ? 1460018 :
    (addr==90) ? 1476465 :
    (addr==91) ? 1492913 :
    (addr==92) ? 1509363 :
    (addr==93) ? 1525814 :
    (addr==94) ? 1542267 :
    (addr==95) ? 1558721 :
    (addr==96) ? 1575177 :
    (addr==97) ? 1591634 :
    (addr==98) ? 1608093 :
    (addr==99) ? 1624553 :
    (addr==100) ? 1641015 :
    (addr==101) ? 1657478 :
    (addr==102) ? 1673943 :
    (addr==103) ? 1690410 :
    (addr==104) ? 1706879 :
    (addr==105) ? 1723349 :
    (addr==106) ? 1739820 :
    (addr==107) ? 1756293 :
    (addr==108) ? 1772769 :
    (addr==109) ? 1789245 :
    (addr==110) ? 1805724 :
    (addr==111) ? 1822204 :
    (addr==112) ? 1838686 :
    (addr==113) ? 1855170 :
    (addr==114) ? 1871655 :
    (addr==115) ? 1888143 :
    (addr==116) ? 1904632 :
    (addr==117) ? 1921123 :
    (addr==118) ? 1937616 :
    (addr==119) ? 1954111 :
    (addr==120) ? 1970608 :
    (addr==121) ? 1987106 :
    (addr==122) ? 2003607 :
    (addr==123) ? 2020109 :
    (addr==124) ? 2036614 :
    (addr==125) ? 2053120 :
    (addr==126) ? 2069629 :
    (addr==127) ? 2086139 :
    (addr==128) ? 2102652 :
    (addr==129) ? 2119166 :
    (addr==130) ? 2135683 :
    (addr==131) ? 2152201 :
    (addr==132) ? 2168722 :
    (addr==133) ? 2185245 :
    (addr==134) ? 2201770 :
    (addr==135) ? 2218297 :
    (addr==136) ? 2234827 :
    (addr==137) ? 2251358 :
    (addr==138) ? 2267892 :
    (addr==139) ? 2284428 :
    (addr==140) ? 2300966 :
    (addr==141) ? 2317507 :
    (addr==142) ? 2334049 :
    (addr==143) ? 2350594 :
    (addr==144) ? 2367142 :
    (addr==145) ? 2383691 :
    (addr==146) ? 2400243 :
    (addr==147) ? 2416797 :
    (addr==148) ? 2433354 :
    (addr==149) ? 2449913 :
    (addr==150) ? 2466475 :
    (addr==151) ? 2483038 :
    (addr==152) ? 2499605 :
    (addr==153) ? 2516173 :
    (addr==154) ? 2532745 :
    (addr==155) ? 2549318 :
    (addr==156) ? 2565895 :
    (addr==157) ? 2582473 :
    (addr==158) ? 2599055 :
    (addr==159) ? 2615639 :
    (addr==160) ? 2632225 :
    (addr==161) ? 2648814 :
    (addr==162) ? 2665406 :
    (addr==163) ? 2682000 :
    (addr==164) ? 2698597 :
    (addr==165) ? 2715197 :
    (addr==166) ? 2731799 :
    (addr==167) ? 2748404 :
    (addr==168) ? 2765012 :
    (addr==169) ? 2781622 :
    (addr==170) ? 2798235 :
    (addr==171) ? 2814851 :
    (addr==172) ? 2831470 :
    (addr==173) ? 2848091 :
    (addr==174) ? 2864716 :
    (addr==175) ? 2881343 :
    (addr==176) ? 2897973 :
    (addr==177) ? 2914606 :
    (addr==178) ? 2931242 :
    (addr==179) ? 2947880 :
    (addr==180) ? 2964522 :
    (addr==181) ? 2981167 :
    (addr==182) ? 2997814 :
    (addr==183) ? 3014465 :
    (addr==184) ? 3031119 :
    (addr==185) ? 3047775 :
    (addr==186) ? 3064435 :
    (addr==187) ? 3081097 :
    (addr==188) ? 3097763 :
    (addr==189) ? 3114432 :
    (addr==190) ? 3131104 :
    (addr==191) ? 3147779 :
    (addr==192) ? 3164457 :
    (addr==193) ? 3181139 :
    (addr==194) ? 3197823 :
    (addr==195) ? 3214511 :
    (addr==196) ? 3231202 :
    (addr==197) ? 3247896 :
    (addr==198) ? 3264594 :
    (addr==199) ? 3281295 :
    (addr==200) ? 3297999 :
    (addr==201) ? 3314706 :
    (addr==202) ? 3331417 :
    (addr==203) ? 3348131 :
    (addr==204) ? 3364848 :
    (addr==205) ? 3381569 :
    (addr==206) ? 3398294 :
    (addr==207) ? 3415021 :
    (addr==208) ? 3431752 :
    (addr==209) ? 3448487 :
    (addr==210) ? 3465225 :
    (addr==211) ? 3481966 :
    (addr==212) ? 3498711 :
    (addr==213) ? 3515460 :
    (addr==214) ? 3532212 :
    (addr==215) ? 3548968 :
    (addr==216) ? 3565727 :
    (addr==217) ? 3582490 :
    (addr==218) ? 3599257 :
    (addr==219) ? 3616027 :
    (addr==220) ? 3632801 :
    (addr==221) ? 3649579 :
    (addr==222) ? 3666360 :
    (addr==223) ? 3683145 :
    (addr==224) ? 3699934 :
    (addr==225) ? 3716726 :
    (addr==226) ? 3733523 :
    (addr==227) ? 3750323 :
    (addr==228) ? 3767127 :
    (addr==229) ? 3783934 :
    (addr==230) ? 3800746 :
    (addr==231) ? 3817562 :
    (addr==232) ? 3834381 :
    (addr==233) ? 3851204 :
    (addr==234) ? 3868032 :
    (addr==235) ? 3884863 :
    (addr==236) ? 3901698 :
    (addr==237) ? 3918538 :
    (addr==238) ? 3935381 :
    (addr==239) ? 3952228 :
    (addr==240) ? 3969080 :
    (addr==241) ? 3985935 :
    (addr==242) ? 4002795 :
    (addr==243) ? 4019658 :
    (addr==244) ? 4036526 :
    (addr==245) ? 4053398 :
    (addr==246) ? 4070274 :
    (addr==247) ? 4087155 :
    (addr==248) ? 4104039 :
    (addr==249) ? 4120928 :
    (addr==250) ? 4137821 :
    (addr==251) ? 4154719 :
    (addr==252) ? 4171620 :
    (addr==253) ? 4188526 :
    (addr==254) ? 4205437 :
    (addr==255) ? 4222352 :
    (addr==256) ? 4239271 :
    (addr==257) ? 4256194 :
    (addr==258) ? 4273122 :
    (addr==259) ? 4290055 :
    (addr==260) ? 4306991 :
    (addr==261) ? 4323933 :
    (addr==262) ? 4340879 :
    (addr==263) ? 4357829 :
    (addr==264) ? 4374784 :
    (addr==265) ? 4391744 :
    (addr==266) ? 4408708 :
    (addr==267) ? 4425676 :
    (addr==268) ? 4442650 :
    (addr==269) ? 4459628 :
    (addr==270) ? 4476611 :
    (addr==271) ? 4493598 :
    (addr==272) ? 4510590 :
    (addr==273) ? 4527587 :
    (addr==274) ? 4544589 :
    (addr==275) ? 4561595 :
    (addr==276) ? 4578606 :
    (addr==277) ? 4595622 :
    (addr==278) ? 4612643 :
    (addr==279) ? 4629669 :
    (addr==280) ? 4646700 :
    (addr==281) ? 4663735 :
    (addr==282) ? 4680776 :
    (addr==283) ? 4697821 :
    (addr==284) ? 4714872 :
    (addr==285) ? 4731927 :
    (addr==286) ? 4748988 :
    (addr==287) ? 4766053 :
    (addr==288) ? 4783124 :
    (addr==289) ? 4800200 :
    (addr==290) ? 4817281 :
    (addr==291) ? 4834367 :
    (addr==292) ? 4851458 :
    (addr==293) ? 4868554 :
    (addr==294) ? 4885656 :
    (addr==295) ? 4902762 :
    (addr==296) ? 4919874 :
    (addr==297) ? 4936992 :
    (addr==298) ? 4954114 :
    (addr==299) ? 4971242 :
    (addr==300) ? 4988375 :
    (addr==301) ? 5005514 :
    (addr==302) ? 5022658 :
    (addr==303) ? 5039807 :
    (addr==304) ? 5056962 :
    (addr==305) ? 5074122 :
    (addr==306) ? 5091288 :
    (addr==307) ? 5108459 :
    (addr==308) ? 5125636 :
    (addr==309) ? 5142818 :
    (addr==310) ? 5160006 :
    (addr==311) ? 5177199 :
    (addr==312) ? 5194399 :
    (addr==313) ? 5211603 :
    (addr==314) ? 5228814 :
    (addr==315) ? 5246030 :
    (addr==316) ? 5263252 :
    (addr==317) ? 5280479 :
    (addr==318) ? 5297712 :
    (addr==319) ? 5314952 :
    (addr==320) ? 5332196 :
    (addr==321) ? 5349447 :
    (addr==322) ? 5366704 :
    (addr==323) ? 5383966 :
    (addr==324) ? 5401235 :
    (addr==325) ? 5418509 :
    (addr==326) ? 5435789 :
    (addr==327) ? 5453075 :
    (addr==328) ? 5470368 :
    (addr==329) ? 5487666 :
    (addr==330) ? 5504970 :
    (addr==331) ? 5522281 :
    (addr==332) ? 5539597 :
    (addr==333) ? 5556920 :
    (addr==334) ? 5574249 :
    (addr==335) ? 5591584 :
    (addr==336) ? 5608925 :
    (addr==337) ? 5626272 :
    (addr==338) ? 5643626 :
    (addr==339) ? 5660986 :
    (addr==340) ? 5678352 :
    (addr==341) ? 5695724 :
    (addr==342) ? 5713103 :
    (addr==343) ? 5730489 :
    (addr==344) ? 5747880 :
    (addr==345) ? 5765279 :
    (addr==346) ? 5782683 :
    (addr==347) ? 5800094 :
    (addr==348) ? 5817512 :
    (addr==349) ? 5834936 :
    (addr==350) ? 5852367 :
    (addr==351) ? 5869804 :
    (addr==352) ? 5887248 :
    (addr==353) ? 5904698 :
    (addr==354) ? 5922156 :
    (addr==355) ? 5939619 :
    (addr==356) ? 5957090 :
    (addr==357) ? 5974567 :
    (addr==358) ? 5992052 :
    (addr==359) ? 6009543 :
    (addr==360) ? 6027040 :
    (addr==361) ? 6044545 :
    (addr==362) ? 6062056 :
    (addr==363) ? 6079575 :
    (addr==364) ? 6097100 :
    (addr==365) ? 6114633 :
    (addr==366) ? 6132172 :
    (addr==367) ? 6149718 :
    (addr==368) ? 6167272 :
    (addr==369) ? 6184832 :
    (addr==370) ? 6202400 :
    (addr==371) ? 6219974 :
    (addr==372) ? 6237556 :
    (addr==373) ? 6255145 :
    (addr==374) ? 6272742 :
    (addr==375) ? 6290345 :
    (addr==376) ? 6307956 :
    (addr==377) ? 6325574 :
    (addr==378) ? 6343199 :
    (addr==379) ? 6360832 :
    (addr==380) ? 6378472 :
    (addr==381) ? 6396120 :
    (addr==382) ? 6413775 :
    (addr==383) ? 6431437 :
    (addr==384) ? 6449107 :
    (addr==385) ? 6466785 :
    (addr==386) ? 6484470 :
    (addr==387) ? 6502162 :
    (addr==388) ? 6519863 :
    (addr==389) ? 6537571 :
    (addr==390) ? 6555286 :
    (addr==391) ? 6573010 :
    (addr==392) ? 6590741 :
    (addr==393) ? 6608480 :
    (addr==394) ? 6626226 :
    (addr==395) ? 6643981 :
    (addr==396) ? 6661743 :
    (addr==397) ? 6679513 :
    (addr==398) ? 6697291 :
    (addr==399) ? 6715077 :
    (addr==400) ? 6732871 :
    (addr==401) ? 6750673 :
    (addr==402) ? 6768484 :
    (addr==403) ? 6786302 :
    (addr==404) ? 6804128 :
    (addr==405) ? 6821962 :
    (addr==406) ? 6839805 :
    (addr==407) ? 6857656 :
    (addr==408) ? 6875515 :
    (addr==409) ? 6893382 :
    (addr==410) ? 6911258 :
    (addr==411) ? 6929142 :
    (addr==412) ? 6947034 :
    (addr==413) ? 6964935 :
    (addr==414) ? 6982844 :
    (addr==415) ? 7000761 :
    (addr==416) ? 7018687 :
    (addr==417) ? 7036622 :
    (addr==418) ? 7054565 :
    (addr==419) ? 7072516 :
    (addr==420) ? 7090477 :
    (addr==421) ? 7108446 :
    (addr==422) ? 7126423 :
    (addr==423) ? 7144410 :
    (addr==424) ? 7162405 :
    (addr==425) ? 7180409 :
    (addr==426) ? 7198421 :
    (addr==427) ? 7216443 :
    (addr==428) ? 7234473 :
    (addr==429) ? 7252513 :
    (addr==430) ? 7270561 :
    (addr==431) ? 7288618 :
    (addr==432) ? 7306685 :
    (addr==433) ? 7324760 :
    (addr==434) ? 7342844 :
    (addr==435) ? 7360938 :
    (addr==436) ? 7379041 :
    (addr==437) ? 7397153 :
    (addr==438) ? 7415274 :
    (addr==439) ? 7433404 :
    (addr==440) ? 7451544 :
    (addr==441) ? 7469693 :
    (addr==442) ? 7487852 :
    (addr==443) ? 7506020 :
    (addr==444) ? 7524197 :
    (addr==445) ? 7542384 :
    (addr==446) ? 7560580 :
    (addr==447) ? 7578786 :
    (addr==448) ? 7597001 :
    (addr==449) ? 7615226 :
    (addr==450) ? 7633461 :
    (addr==451) ? 7651706 :
    (addr==452) ? 7669960 :
    (addr==453) ? 7688224 :
    (addr==454) ? 7706498 :
    (addr==455) ? 7724781 :
    (addr==456) ? 7743075 :
    (addr==457) ? 7761378 :
    (addr==458) ? 7779692 :
    (addr==459) ? 7798015 :
    (addr==460) ? 7816348 :
    (addr==461) ? 7834692 :
    (addr==462) ? 7853046 :
    (addr==463) ? 7871409 :
    (addr==464) ? 7889783 :
    (addr==465) ? 7908168 :
    (addr==466) ? 7926562 :
    (addr==467) ? 7944967 :
    (addr==468) ? 7963382 :
    (addr==469) ? 7981808 :
    (addr==470) ? 8000244 :
    (addr==471) ? 8018690 :
    (addr==472) ? 8037147 :
    (addr==473) ? 8055615 :
    (addr==474) ? 8074093 :
    (addr==475) ? 8092582 :
    (addr==476) ? 8111081 :
    (addr==477) ? 8129591 :
    (addr==478) ? 8148112 :
    (addr==479) ? 8166644 :
    (addr==480) ? 8185186 :
    (addr==481) ? 8203740 :
    (addr==482) ? 8222304 :
    (addr==483) ? 8240879 :
    (addr==484) ? 8259466 :
    (addr==485) ? 8278063 :
    (addr==486) ? 8296671 :
    (addr==487) ? 8315291 :
    (addr==488) ? 8333922 :
    (addr==489) ? 8352564 :
    (addr==490) ? 8371217 :
    (addr==491) ? 8389882 :
    (addr==492) ? 8408558 :
    (addr==493) ? 8427245 :
    (addr==494) ? 8445944 :
    (addr==495) ? 8464654 :
    (addr==496) ? 8483376 :
    (addr==497) ? 8502109 :
    (addr==498) ? 8520854 :
    (addr==499) ? 8539611 :
    (addr==500) ? 8558379 :
    (addr==501) ? 8577159 :
    (addr==502) ? 8595951 :
    (addr==503) ? 8614755 :
    (addr==504) ? 8633570 :
    (addr==505) ? 8652398 :
    (addr==506) ? 8671238 :
    (addr==507) ? 8690089 :
    (addr==508) ? 8708953 :
    (addr==509) ? 8727829 :
    (addr==510) ? 8746717 :
    (addr==511) ? 8765617 :
    (addr==512) ? 8784529 :
    (addr==513) ? 8803454 :
    (addr==514) ? 8822391 :
    (addr==515) ? 8841341 :
    (addr==516) ? 8860303 :
    (addr==517) ? 8879277 :
    (addr==518) ? 8898264 :
    (addr==519) ? 8917264 :
    (addr==520) ? 8936276 :
    (addr==521) ? 8955302 :
    (addr==522) ? 8974339 :
    (addr==523) ? 8993390 :
    (addr==524) ? 9012453 :
    (addr==525) ? 9031530 :
    (addr==526) ? 9050619 :
    (addr==527) ? 9069722 :
    (addr==528) ? 9088837 :
    (addr==529) ? 9107966 :
    (addr==530) ? 9127107 :
    (addr==531) ? 9146262 :
    (addr==532) ? 9165431 :
    (addr==533) ? 9184612 :
    (addr==534) ? 9203807 :
    (addr==535) ? 9223015 :
    (addr==536) ? 9242237 :
    (addr==537) ? 9261473 :
    (addr==538) ? 9280722 :
    (addr==539) ? 9299984 :
    (addr==540) ? 9319260 :
    (addr==541) ? 9338551 :
    (addr==542) ? 9357854 :
    (addr==543) ? 9377172 :
    (addr==544) ? 9396504 :
    (addr==545) ? 9415850 :
    (addr==546) ? 9435209 :
    (addr==547) ? 9454583 :
    (addr==548) ? 9473971 :
    (addr==549) ? 9493373 :
    (addr==550) ? 9512789 :
    (addr==551) ? 9532220 :
    (addr==552) ? 9551665 :
    (addr==553) ? 9571125 :
    (addr==554) ? 9590599 :
    (addr==555) ? 9610087 :
    (addr==556) ? 9629591 :
    (addr==557) ? 9649108 :
    (addr==558) ? 9668641 :
    (addr==559) ? 9688188 :
    (addr==560) ? 9707751 :
    (addr==561) ? 9727328 :
    (addr==562) ? 9746920 :
    (addr==563) ? 9766527 :
    (addr==564) ? 9786149 :
    (addr==565) ? 9805786 :
    (addr==566) ? 9825439 :
    (addr==567) ? 9845107 :
    (addr==568) ? 9864790 :
    (addr==569) ? 9884489 :
    (addr==570) ? 9904203 :
    (addr==571) ? 9923933 :
    (addr==572) ? 9943678 :
    (addr==573) ? 9963439 :
    (addr==574) ? 9983215 :
    (addr==575) ? 10003008 :
    (addr==576) ? 10022816 :
    (addr==577) ? 10042640 :
    (addr==578) ? 10062480 :
    (addr==579) ? 10082337 :
    (addr==580) ? 10102209 :
    (addr==581) ? 10122098 :
    (addr==582) ? 10142002 :
    (addr==583) ? 10161924 :
    (addr==584) ? 10181861 :
    (addr==585) ? 10201815 :
    (addr==586) ? 10221786 :
    (addr==587) ? 10241773 :
    (addr==588) ? 10261777 :
    (addr==589) ? 10281797 :
    (addr==590) ? 10301834 :
    (addr==591) ? 10321889 :
    (addr==592) ? 10341960 :
    (addr==593) ? 10362048 :
    (addr==594) ? 10382153 :
    (addr==595) ? 10402276 :
    (addr==596) ? 10422416 :
    (addr==597) ? 10442573 :
    (addr==598) ? 10462747 :
    (addr==599) ? 10482939 :
    (addr==600) ? 10503149 :
    (addr==601) ? 10523376 :
    (addr==602) ? 10543621 :
    (addr==603) ? 10563883 :
    (addr==604) ? 10584163 :
    (addr==605) ? 10604462 :
    (addr==606) ? 10624778 :
    (addr==607) ? 10645112 :
    (addr==608) ? 10665465 :
    (addr==609) ? 10685836 :
    (addr==610) ? 10706225 :
    (addr==611) ? 10726632 :
    (addr==612) ? 10747058 :
    (addr==613) ? 10767503 :
    (addr==614) ? 10787966 :
    (addr==615) ? 10808448 :
    (addr==616) ? 10828949 :
    (addr==617) ? 10849468 :
    (addr==618) ? 10870007 :
    (addr==619) ? 10890564 :
    (addr==620) ? 10911141 :
    (addr==621) ? 10931737 :
    (addr==622) ? 10952352 :
    (addr==623) ? 10972987 :
    (addr==624) ? 10993641 :
    (addr==625) ? 11014315 :
    (addr==626) ? 11035008 :
    (addr==627) ? 11055721 :
    (addr==628) ? 11076454 :
    (addr==629) ? 11097206 :
    (addr==630) ? 11117979 :
    (addr==631) ? 11138772 :
    (addr==632) ? 11159585 :
    (addr==633) ? 11180418 :
    (addr==634) ? 11201272 :
    (addr==635) ? 11222146 :
    (addr==636) ? 11243041 :
    (addr==637) ? 11263956 :
    (addr==638) ? 11284892 :
    (addr==639) ? 11305849 :
    (addr==640) ? 11326827 :
    (addr==641) ? 11347826 :
    (addr==642) ? 11368846 :
    (addr==643) ? 11389887 :
    (addr==644) ? 11410950 :
    (addr==645) ? 11432033 :
    (addr==646) ? 11453139 :
    (addr==647) ? 11474266 :
    (addr==648) ? 11495415 :
    (addr==649) ? 11516585 :
    (addr==650) ? 11537778 :
    (addr==651) ? 11558992 :
    (addr==652) ? 11580229 :
    (addr==653) ? 11601487 :
    (addr==654) ? 11622769 :
    (addr==655) ? 11644072 :
    (addr==656) ? 11665398 :
    (addr==657) ? 11686747 :
    (addr==658) ? 11708118 :
    (addr==659) ? 11729513 :
    (addr==660) ? 11750930 :
    (addr==661) ? 11772370 :
    (addr==662) ? 11793834 :
    (addr==663) ? 11815321 :
    (addr==664) ? 11836831 :
    (addr==665) ? 11858365 :
    (addr==666) ? 11879922 :
    (addr==667) ? 11901503 :
    (addr==668) ? 11923108 :
    (addr==669) ? 11944737 :
    (addr==670) ? 11966390 :
    (addr==671) ? 11988068 :
    (addr==672) ? 12009769 :
    (addr==673) ? 12031495 :
    (addr==674) ? 12053246 :
    (addr==675) ? 12075021 :
    (addr==676) ? 12096821 :
    (addr==677) ? 12118646 :
    (addr==678) ? 12140496 :
    (addr==679) ? 12162372 :
    (addr==680) ? 12184272 :
    (addr==681) ? 12206198 :
    (addr==682) ? 12228149 :
    (addr==683) ? 12250127 :
    (addr==684) ? 12272130 :
    (addr==685) ? 12294158 :
    (addr==686) ? 12316213 :
    (addr==687) ? 12338295 :
    (addr==688) ? 12360402 :
    (addr==689) ? 12382536 :
    (addr==690) ? 12404696 :
    (addr==691) ? 12426884 :
    (addr==692) ? 12449098 :
    (addr==693) ? 12471339 :
    (addr==694) ? 12493607 :
    (addr==695) ? 12515903 :
    (addr==696) ? 12538226 :
    (addr==697) ? 12560576 :
    (addr==698) ? 12582954 :
    (addr==699) ? 12605360 :
    (addr==700) ? 12627794 :
    (addr==701) ? 12650256 :
    (addr==702) ? 12672747 :
    (addr==703) ? 12695266 :
    (addr==704) ? 12717813 :
    (addr==705) ? 12740389 :
    (addr==706) ? 12762994 :
    (addr==707) ? 12785628 :
    (addr==708) ? 12808292 :
    (addr==709) ? 12830984 :
    (addr==710) ? 12853706 :
    (addr==711) ? 12876458 :
    (addr==712) ? 12899239 :
    (addr==713) ? 12922051 :
    (addr==714) ? 12944893 :
    (addr==715) ? 12967765 :
    (addr==716) ? 12990667 :
    (addr==717) ? 13013600 :
    (addr==718) ? 13036564 :
    (addr==719) ? 13059558 :
    (addr==720) ? 13082584 :
    (addr==721) ? 13105641 :
    (addr==722) ? 13128730 :
    (addr==723) ? 13151850 :
    (addr==724) ? 13175002 :
    (addr==725) ? 13198186 :
    (addr==726) ? 13221402 :
    (addr==727) ? 13244651 :
    (addr==728) ? 13267932 :
    (addr==729) ? 13291246 :
    (addr==730) ? 13314592 :
    (addr==731) ? 13337972 :
    (addr==732) ? 13361385 :
    (addr==733) ? 13384831 :
    (addr==734) ? 13408312 :
    (addr==735) ? 13431825 :
    (addr==736) ? 13455373 :
    (addr==737) ? 13478955 :
    (addr==738) ? 13502572 :
    (addr==739) ? 13526223 :
    (addr==740) ? 13549909 :
    (addr==741) ? 13573630 :
    (addr==742) ? 13597386 :
    (addr==743) ? 13621178 :
    (addr==744) ? 13645005 :
    (addr==745) ? 13668868 :
    (addr==746) ? 13692767 :
    (addr==747) ? 13716703 :
    (addr==748) ? 13740675 :
    (addr==749) ? 13764683 :
    (addr==750) ? 13788729 :
    (addr==751) ? 13812811 :
    (addr==752) ? 13836931 :
    (addr==753) ? 13861089 :
    (addr==754) ? 13885284 :
    (addr==755) ? 13909518 :
    (addr==756) ? 13933789 :
    (addr==757) ? 13958099 :
    (addr==758) ? 13982448 :
    (addr==759) ? 14006836 :
    (addr==760) ? 14031263 :
    (addr==761) ? 14055729 :
    (addr==762) ? 14080236 :
    (addr==763) ? 14104782 :
    (addr==764) ? 14129368 :
    (addr==765) ? 14153995 :
    (addr==766) ? 14178662 :
    (addr==767) ? 14203371 :
    (addr==768) ? 14228120 :
    (addr==769) ? 14252911 :
    (addr==770) ? 14277744 :
    (addr==771) ? 14302619 :
    (addr==772) ? 14327536 :
    (addr==773) ? 14352495 :
    (addr==774) ? 14377498 :
    (addr==775) ? 14402543 :
    (addr==776) ? 14427632 :
    (addr==777) ? 14452765 :
    (addr==778) ? 14477941 :
    (addr==779) ? 14503162 :
    (addr==780) ? 14528427 :
    (addr==781) ? 14553737 :
    (addr==782) ? 14579092 :
    (addr==783) ? 14604493 :
    (addr==784) ? 14629939 :
    (addr==785) ? 14655431 :
    (addr==786) ? 14680970 :
    (addr==787) ? 14706555 :
    (addr==788) ? 14732187 :
    (addr==789) ? 14757867 :
    (addr==790) ? 14783594 :
    (addr==791) ? 14809369 :
    (addr==792) ? 14835192 :
    (addr==793) ? 14861064 :
    (addr==794) ? 14886984 :
    (addr==795) ? 14912954 :
    (addr==796) ? 14938974 :
    (addr==797) ? 14965044 :
    (addr==798) ? 14991163 :
    (addr==799) ? 15017334 :
    (addr==800) ? 15043556 :
    (addr==801) ? 15069829 :
    (addr==802) ? 15096153 :
    (addr==803) ? 15122530 :
    (addr==804) ? 15148960 :
    (addr==805) ? 15175442 :
    (addr==806) ? 15201977 :
    (addr==807) ? 15228567 :
    (addr==808) ? 15255210 :
    (addr==809) ? 15281908 :
    (addr==810) ? 15308660 :
    (addr==811) ? 15335468 :
    (addr==812) ? 15362332 :
    (addr==813) ? 15389251 :
    (addr==814) ? 15416228 :
    (addr==815) ? 15443261 :
    (addr==816) ? 15470351 :
    (addr==817) ? 15497500 :
    (addr==818) ? 15524706 :
    (addr==819) ? 15551972 :
    (addr==820) ? 15579296 :
    (addr==821) ? 15606680 :
    (addr==822) ? 15634124 :
    (addr==823) ? 15661629 :
    (addr==824) ? 15689195 :
    (addr==825) ? 15716822 :
    (addr==826) ? 15744512 :
    (addr==827) ? 15772263 :
    (addr==828) ? 15800078 :
    (addr==829) ? 15827957 :
    (addr==830) ? 15855899 :
    (addr==831) ? 15883906 :
    (addr==832) ? 15911978 :
    (addr==833) ? 15940116 :
    (addr==834) ? 15968320 :
    (addr==835) ? 15996590 :
    (addr==836) ? 16024928 :
    (addr==837) ? 16053334 :
    (addr==838) ? 16081808 :
    (addr==839) ? 16110351 :
    (addr==840) ? 16138963 :
    (addr==841) ? 16167646 :
    (addr==842) ? 16196400 :
    (addr==843) ? 16225225 :
    (addr==844) ? 16254122 :
    (addr==845) ? 16283091 :
    (addr==846) ? 16312134 :
    (addr==847) ? 16341251 :
    (addr==848) ? 16370442 :
    (addr==849) ? 16399708 :
    (addr==850) ? 16429051 :
    (addr==851) ? 16458470 :
    (addr==852) ? 16487966 :
    (addr==853) ? 16517540 :
    (addr==854) ? 16547193 :
    (addr==855) ? 16576926 :
    (addr==856) ? 16606738 :
    (addr==857) ? 16636632 :
    (addr==858) ? 16666607 :
    (addr==859) ? 16696664 :
    (addr==860) ? 16726805 :
    (addr==861) ? 16757030 :
    (addr==862) ? 16787340 :
    (addr==863) ? 16817735 :
    (addr==864) ? 16848217 :
    (addr==865) ? 16878786 :
    (addr==866) ? 16909443 :
    (addr==867) ? 16940189 :
    (addr==868) ? 16971025 :
    (addr==869) ? 17001952 :
    (addr==870) ? 17032971 :
    (addr==871) ? 17064082 :
    (addr==872) ? 17095287 :
    (addr==873) ? 17126587 :
    (addr==874) ? 17157982 :
    (addr==875) ? 17189473 :
    (addr==876) ? 17221062 :
    (addr==877) ? 17252750 :
    (addr==878) ? 17284537 :
    (addr==879) ? 17316425 :
    (addr==880) ? 17348415 :
    (addr==881) ? 17380508 :
    (addr==882) ? 17412704 :
    (addr==883) ? 17445006 :
    (addr==884) ? 17477414 :
    (addr==885) ? 17509929 :
    (addr==886) ? 17542553 :
    (addr==887) ? 17575286 :
    (addr==888) ? 17608131 :
    (addr==889) ? 17641089 :
    (addr==890) ? 17674159 :
    (addr==891) ? 17707345 :
    (addr==892) ? 17740647 :
    (addr==893) ? 17774067 :
    (addr==894) ? 17807606 :
    (addr==895) ? 17841265 :
    (addr==896) ? 17875046 :
    (addr==897) ? 17908951 :
    (addr==898) ? 17942980 :
    (addr==899) ? 17977136 :
    (addr==900) ? 18011420 :
    (addr==901) ? 18045834 :
    (addr==902) ? 18080378 :
    (addr==903) ? 18115056 :
    (addr==904) ? 18149868 :
    (addr==905) ? 18184816 :
    (addr==906) ? 18219903 :
    (addr==907) ? 18255129 :
    (addr==908) ? 18290497 :
    (addr==909) ? 18326009 :
    (addr==910) ? 18361666 :
    (addr==911) ? 18397470 :
    (addr==912) ? 18433424 :
    (addr==913) ? 18469530 :
    (addr==914) ? 18505789 :
    (addr==915) ? 18542204 :
    (addr==916) ? 18578777 :
    (addr==917) ? 18615511 :
    (addr==918) ? 18652407 :
    (addr==919) ? 18689467 :
    (addr==920) ? 18726695 :
    (addr==921) ? 18764093 :
    (addr==922) ? 18801663 :
    (addr==923) ? 18839409 :
    (addr==924) ? 18877331 :
    (addr==925) ? 18915434 :
    (addr==926) ? 18953720 :
    (addr==927) ? 18992193 :
    (addr==928) ? 19030854 :
    (addr==929) ? 19069707 :
    (addr==930) ? 19108755 :
    (addr==931) ? 19148001 :
    (addr==932) ? 19187448 :
    (addr==933) ? 19227101 :
    (addr==934) ? 19266962 :
    (addr==935) ? 19307034 :
    (addr==936) ? 19347323 :
    (addr==937) ? 19387830 :
    (addr==938) ? 19428561 :
    (addr==939) ? 19469518 :
    (addr==940) ? 19510707 :
    (addr==941) ? 19552131 :
    (addr==942) ? 19593795 :
    (addr==943) ? 19635702 :
    (addr==944) ? 19677859 :
    (addr==945) ? 19720269 :
    (addr==946) ? 19762938 :
    (addr==947) ? 19805870 :
    (addr==948) ? 19849071 :
    (addr==949) ? 19892546 :
    (addr==950) ? 19936301 :
    (addr==951) ? 19980341 :
    (addr==952) ? 20024673 :
    (addr==953) ? 20069302 :
    (addr==954) ? 20114236 :
    (addr==955) ? 20159480 :
    (addr==956) ? 20205042 :
    (addr==957) ? 20250928 :
    (addr==958) ? 20297146 :
    (addr==959) ? 20343705 :
    (addr==960) ? 20390610 :
    (addr==961) ? 20437872 :
    (addr==962) ? 20485499 :
    (addr==963) ? 20533499 :
    (addr==964) ? 20581882 :
    (addr==965) ? 20630657 :
    (addr==966) ? 20679836 :
    (addr==967) ? 20729427 :
    (addr==968) ? 20779443 :
    (addr==969) ? 20829896 :
    (addr==970) ? 20880796 :
    (addr==971) ? 20932156 :
    (addr==972) ? 20983991 :
    (addr==973) ? 21036313 :
    (addr==974) ? 21089138 :
    (addr==975) ? 21142480 :
    (addr==976) ? 21196356 :
    (addr==977) ? 21250782 :
    (addr==978) ? 21305777 :
    (addr==979) ? 21361359 :
    (addr==980) ? 21417548 :
    (addr==981) ? 21474365 :
    (addr==982) ? 21531832 :
    (addr==983) ? 21589974 :
    (addr==984) ? 21648814 :
    (addr==985) ? 21708379 :
    (addr==986) ? 21768698 :
    (addr==987) ? 21829801 :
    (addr==988) ? 21891720 :
    (addr==989) ? 21954489 :
    (addr==990) ? 22018146 :
    (addr==991) ? 22082731 :
    (addr==992) ? 22148285 :
    (addr==993) ? 22214855 :
    (addr==994) ? 22282491 :
    (addr==995) ? 22351247 :
    (addr==996) ? 22421181 :
    (addr==997) ? 22492358 :
    (addr==998) ? 22564849 :
    (addr==999) ? 22638729 :
    (addr==1000) ? 22714083 :
    (addr==1001) ? 22791005 :
    (addr==1002) ? 22869599 :
    (addr==1003) ? 22949980 :
    (addr==1004) ? 23032279 :
    (addr==1005) ? 23116642 :
    (addr==1006) ? 23203234 :
    (addr==1007) ? 23292245 :
    (addr==1008) ? 23383893 :
    (addr==1009) ? 23478428 :
    (addr==1010) ? 23576147 :
    (addr==1011) ? 23677398 :
    (addr==1012) ? 23782598 :
    (addr==1013) ? 23892253 :
    (addr==1014) ? 24006989 :
    (addr==1015) ? 24127591 :
    (addr==1016) ? 24255069 :
    (addr==1017) ? 24390763 :
    (addr==1018) ? 24536514 :
    (addr==1019) ? 24694969 :
    (addr==1020) ? 24870195 :
    (addr==1021) ? 25069037 :
    (addr==1022) ? 25304842 :
    (addr==1023) ? 25612073 :
25'bx;
endmodule
